<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-102.213,106.838,146.413,-153.038</PageViewport>
<gate>
<ID>1</ID>
<type>DA_FROM</type>
<position>68,-28.5</position>
<input>
<ID>IN_0</ID>235 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND2</lparam></gate>
<gate>
<ID>2</ID>
<type>DA_FROM</type>
<position>48.5,56</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>3</ID>
<type>DA_FROM</type>
<position>40,44.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>4</ID>
<type>DA_FROM</type>
<position>73,-16.5</position>
<input>
<ID>IN_0</ID>224 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>5</ID>
<type>DE_TO</type>
<position>80,42.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0</lparam></gate>
<gate>
<ID>6</ID>
<type>DA_FROM</type>
<position>20,17</position>
<input>
<ID>IN_0</ID>64 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>7</ID>
<type>DA_FROM</type>
<position>58,15.5</position>
<input>
<ID>IN_0</ID>218 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>8</ID>
<type>AM_MUX_16x1</type>
<position>74.5,42.5</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>70 </input>
<input>
<ID>IN_10</ID>173 </input>
<input>
<ID>IN_11</ID>202 </input>
<input>
<ID>IN_12</ID>200 </input>
<input>
<ID>IN_13</ID>201 </input>
<input>
<ID>IN_14</ID>199 </input>
<input>
<ID>IN_15</ID>198 </input>
<input>
<ID>IN_2</ID>71 </input>
<input>
<ID>IN_3</ID>72 </input>
<input>
<ID>IN_4</ID>74 </input>
<input>
<ID>IN_5</ID>75 </input>
<input>
<ID>IN_6</ID>98 </input>
<input>
<ID>IN_7</ID>98 </input>
<input>
<ID>IN_8</ID>171 </input>
<input>
<ID>IN_9</ID>172 </input>
<output>
<ID>OUT</ID>1 </output>
<input>
<ID>SEL_0</ID>5 </input>
<input>
<ID>SEL_1</ID>4 </input>
<input>
<ID>SEL_2</ID>2 </input>
<input>
<ID>SEL_3</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>9</ID>
<type>DA_FROM</type>
<position>48.5,54</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>10</ID>
<type>DA_FROM</type>
<position>36,44.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>11</ID>
<type>DA_FROM</type>
<position>68,-24.5</position>
<input>
<ID>IN_0</ID>240 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>12</ID>
<type>DA_FROM</type>
<position>76,55</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>13</ID>
<type>DA_FROM</type>
<position>31,44.5</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>14</ID>
<type>DA_FROM</type>
<position>58.5,-32.5</position>
<input>
<ID>IN_0</ID>232 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum2</lparam></gate>
<gate>
<ID>15</ID>
<type>DA_FROM</type>
<position>75,60</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>74,55</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>17</ID>
<type>DA_FROM</type>
<position>75,-16.5</position>
<input>
<ID>IN_0</ID>227 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>73,60</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>19</ID>
<type>DA_FROM</type>
<position>7,12</position>
<input>
<ID>IN_0</ID>42 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>18,44.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>58.5,-30</position>
<input>
<ID>IN_0</ID>234 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec2</lparam></gate>
<gate>
<ID>22</ID>
<type>DA_FROM</type>
<position>16,44.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>23</ID>
<type>DE_TO</type>
<position>7.5,-2.5</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID UF</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>13,44.5</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>25</ID>
<type>DA_FROM</type>
<position>11,44.5</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>26</ID>
<type>DA_FROM</type>
<position>9,44.5</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>27</ID>
<type>DE_TO</type>
<position>28.5,-2</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff3</lparam></gate>
<gate>
<ID>28</ID>
<type>DA_FROM</type>
<position>7,44.5</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>29</ID>
<type>DA_FROM</type>
<position>11,12</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>30</ID>
<type>DE_TO</type>
<position>34.5,30.5</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum0</lparam></gate>
<gate>
<ID>31</ID>
<type>DE_TO</type>
<position>32.5,30.5</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum1</lparam></gate>
<gate>
<ID>32</ID>
<type>DE_TO</type>
<position>11,-2</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff7</lparam></gate>
<gate>
<ID>33</ID>
<type>DE_TO</type>
<position>30.5,30.5</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum2</lparam></gate>
<gate>
<ID>34</ID>
<type>DE_TO</type>
<position>28.5,30.5</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum3</lparam></gate>
<gate>
<ID>35</ID>
<type>DE_TO</type>
<position>17,30.5</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum4</lparam></gate>
<gate>
<ID>36</ID>
<type>DE_TO</type>
<position>15,30.5</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum5</lparam></gate>
<gate>
<ID>37</ID>
<type>DE_TO</type>
<position>13,30.5</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum6</lparam></gate>
<gate>
<ID>38</ID>
<type>DE_TO</type>
<position>11,30.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum7</lparam></gate>
<gate>
<ID>39</ID>
<type>DE_TO</type>
<position>15,-2</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff5</lparam></gate>
<gate>
<ID>40</ID>
<type>FF_GND</type>
<position>40.5,37</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>41</ID>
<type>DE_TO</type>
<position>7.5,30</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID OV</lparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>5.5,30</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum8</lparam></gate>
<gate>
<ID>43</ID>
<type>DA_FROM</type>
<position>13,12</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>44</ID>
<type>DA_FROM</type>
<position>9,12</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_TO</type>
<position>34.5,-2</position>
<input>
<ID>IN_0</ID>43 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff0</lparam></gate>
<gate>
<ID>46</ID>
<type>DA_FROM</type>
<position>20,44.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>32.5,-2</position>
<input>
<ID>IN_0</ID>44 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff1</lparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>30.5,-2</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff2</lparam></gate>
<gate>
<ID>49</ID>
<type>DE_TO</type>
<position>17,-2</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff4</lparam></gate>
<gate>
<ID>50</ID>
<type>DE_TO</type>
<position>13,-2</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff6</lparam></gate>
<gate>
<ID>51</ID>
<type>DE_TO</type>
<position>5.5,-2.5</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff8</lparam></gate>
<gate>
<ID>52</ID>
<type>AE_FULLADDER_4BIT</type>
<position>31.5,5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>36 </input>
<input>
<ID>IN_2</ID>37 </input>
<input>
<ID>IN_3</ID>38 </input>
<input>
<ID>IN_B_0</ID>56 </input>
<input>
<ID>IN_B_1</ID>54 </input>
<input>
<ID>IN_B_2</ID>55 </input>
<input>
<ID>IN_B_3</ID>53 </input>
<output>
<ID>OUT_0</ID>43 </output>
<output>
<ID>OUT_1</ID>44 </output>
<output>
<ID>OUT_2</ID>45 </output>
<output>
<ID>OUT_3</ID>46 </output>
<input>
<ID>carry_in</ID>69 </input>
<output>
<ID>carry_out</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>53</ID>
<type>AE_FULLADDER_4BIT</type>
<position>14,5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>40 </input>
<input>
<ID>IN_2</ID>41 </input>
<input>
<ID>IN_3</ID>42 </input>
<input>
<ID>IN_B_0</ID>65 </input>
<input>
<ID>IN_B_1</ID>66 </input>
<input>
<ID>IN_B_2</ID>67 </input>
<input>
<ID>IN_B_3</ID>68 </input>
<output>
<ID>OUT_0</ID>47 </output>
<output>
<ID>OUT_1</ID>48 </output>
<output>
<ID>OUT_2</ID>49 </output>
<output>
<ID>OUT_3</ID>50 </output>
<input>
<ID>carry_in</ID>34 </input>
<output>
<ID>carry_out</ID>52 </output>
<output>
<ID>overflow</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>54</ID>
<type>DA_FROM</type>
<position>39.5,17</position>
<input>
<ID>IN_0</ID>59 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>55</ID>
<type>DA_FROM</type>
<position>37.5,17</position>
<input>
<ID>IN_0</ID>60 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>56</ID>
<type>DA_FROM</type>
<position>35.5,17</position>
<input>
<ID>IN_0</ID>58 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>57</ID>
<type>DA_FROM</type>
<position>33.5,17</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>31,12</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>59</ID>
<type>DA_FROM</type>
<position>29,12</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>60</ID>
<type>DA_FROM</type>
<position>27,12</position>
<input>
<ID>IN_0</ID>37 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>61</ID>
<type>DA_FROM</type>
<position>25,12</position>
<input>
<ID>IN_0</ID>38 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>62</ID>
<type>AI_INVERTER_4BIT</type>
<position>35,11.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>60 </input>
<input>
<ID>IN_3</ID>59 </input>
<output>
<ID>OUT_0</ID>53 </output>
<output>
<ID>OUT_1</ID>55 </output>
<output>
<ID>OUT_2</ID>54 </output>
<output>
<ID>OUT_3</ID>56 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>63</ID>
<type>DA_FROM</type>
<position>22,17</position>
<input>
<ID>IN_0</ID>63 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>18,17</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>65</ID>
<type>DA_FROM</type>
<position>16,17</position>
<input>
<ID>IN_0</ID>61 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>66</ID>
<type>AI_INVERTER_4BIT</type>
<position>17.5,11.5</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>62 </input>
<input>
<ID>IN_2</ID>64 </input>
<input>
<ID>IN_3</ID>63 </input>
<output>
<ID>OUT_0</ID>68 </output>
<output>
<ID>OUT_1</ID>67 </output>
<output>
<ID>OUT_2</ID>66 </output>
<output>
<ID>OUT_3</ID>65 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>67</ID>
<type>EE_VDD</type>
<position>40.5,8</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>14,56.5</position>
<gparam>LABEL_TEXT ALU</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AE_FULLADDER_4BIT</type>
<position>31.5,37.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>12 </input>
<input>
<ID>IN_2</ID>13 </input>
<input>
<ID>IN_3</ID>14 </input>
<input>
<ID>IN_B_0</ID>7 </input>
<input>
<ID>IN_B_1</ID>8 </input>
<input>
<ID>IN_B_2</ID>9 </input>
<input>
<ID>IN_B_3</ID>10 </input>
<output>
<ID>OUT_0</ID>23 </output>
<output>
<ID>OUT_1</ID>24 </output>
<output>
<ID>OUT_2</ID>25 </output>
<output>
<ID>OUT_3</ID>26 </output>
<input>
<ID>carry_in</ID>31 </input>
<output>
<ID>carry_out</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>70</ID>
<type>AE_FULLADDER_4BIT</type>
<position>14,37.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<input>
<ID>IN_2</ID>21 </input>
<input>
<ID>IN_3</ID>22 </input>
<input>
<ID>IN_B_0</ID>15 </input>
<input>
<ID>IN_B_1</ID>16 </input>
<input>
<ID>IN_B_2</ID>17 </input>
<input>
<ID>IN_B_3</ID>18 </input>
<output>
<ID>OUT_0</ID>27 </output>
<output>
<ID>OUT_1</ID>28 </output>
<output>
<ID>OUT_2</ID>29 </output>
<output>
<ID>OUT_3</ID>30 </output>
<input>
<ID>carry_in</ID>6 </input>
<output>
<ID>carry_out</ID>33 </output>
<output>
<ID>overflow</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>38,44.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>72</ID>
<type>DA_FROM</type>
<position>33.5,44.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>73</ID>
<type>DA_FROM</type>
<position>29,44.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>74</ID>
<type>DA_FROM</type>
<position>27,44.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>75</ID>
<type>DA_FROM</type>
<position>25,44.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>76</ID>
<type>DA_FROM</type>
<position>22,44.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>77</ID>
<type>DE_TO</type>
<position>-14.5,-12.5</position>
<input>
<ID>IN_0</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR5</lparam></gate>
<gate>
<ID>78</ID>
<type>AE_SMALL_INVERTER</type>
<position>63.5,37</position>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>79</ID>
<type>AE_SMALL_INVERTER</type>
<position>68,38</position>
<input>
<ID>IN_0</ID>73 </input>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>-24.5,-39.5</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>81</ID>
<type>DA_FROM</type>
<position>59.5,39</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum0</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>-24.5,-29.5</position>
<input>
<ID>IN_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>49,40</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff0</lparam></gate>
<gate>
<ID>84</ID>
<type>DA_FROM</type>
<position>-24.5,-35.5</position>
<input>
<ID>IN_0</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>85</ID>
<type>DA_FROM</type>
<position>31,-19</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>86</ID>
<type>DA_FROM</type>
<position>13,-19</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>87</ID>
<type>DA_FROM</type>
<position>-24.5,-47.5</position>
<input>
<ID>IN_0</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>88</ID>
<type>DA_FROM</type>
<position>11,-19</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>9,-19</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>90</ID>
<type>DA_FROM</type>
<position>-24.5,-49.5</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>91</ID>
<type>DA_FROM</type>
<position>7,-19</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>92</ID>
<type>DE_TO</type>
<position>33,-43</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec0</lparam></gate>
<gate>
<ID>93</ID>
<type>FF_GND</type>
<position>40.5,-26</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>94</ID>
<type>DE_TO</type>
<position>4.5,-33</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDecOV</lparam></gate>
<gate>
<ID>95</ID>
<type>AE_FULLADDER_4BIT</type>
<position>31.5,-26</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>78 </input>
<input>
<ID>IN_2</ID>79 </input>
<input>
<ID>IN_3</ID>80 </input>
<input>
<ID>IN_B_0</ID>88 </input>
<input>
<ID>IN_B_1</ID>90 </input>
<input>
<ID>IN_B_2</ID>90 </input>
<input>
<ID>IN_B_3</ID>90 </input>
<output>
<ID>OUT_0</ID>85 </output>
<output>
<ID>OUT_1</ID>91 </output>
<output>
<ID>OUT_2</ID>92 </output>
<output>
<ID>OUT_3</ID>93 </output>
<input>
<ID>carry_in</ID>86 </input>
<output>
<ID>carry_out</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>96</ID>
<type>AE_FULLADDER_4BIT</type>
<position>14,-26</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>83 </input>
<input>
<ID>IN_3</ID>84 </input>
<input>
<ID>IN_B_0</ID>89 </input>
<input>
<ID>IN_B_1</ID>89 </input>
<output>
<ID>OUT_0</ID>94 </output>
<output>
<ID>OUT_1</ID>95 </output>
<output>
<ID>OUT_2</ID>96 </output>
<output>
<ID>OUT_3</ID>97 </output>
<input>
<ID>carry_in</ID>76 </input>
<output>
<ID>overflow</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>97</ID>
<type>DA_FROM</type>
<position>29,-19</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>98</ID>
<type>DA_FROM</type>
<position>27,-19</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>99</ID>
<type>DA_FROM</type>
<position>25,-19</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>100</ID>
<type>EE_VDD</type>
<position>37.5,-20</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>101</ID>
<type>DA_FROM</type>
<position>18,-19</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>102</ID>
<type>DA_FROM</type>
<position>33.5,-19</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>103</ID>
<type>DE_TO</type>
<position>32,-32</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec1</lparam></gate>
<gate>
<ID>104</ID>
<type>DE_TO</type>
<position>31,-43</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec2</lparam></gate>
<gate>
<ID>105</ID>
<type>DE_TO</type>
<position>30,-32</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec3</lparam></gate>
<gate>
<ID>106</ID>
<type>DE_TO</type>
<position>15.5,-32</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec4</lparam></gate>
<gate>
<ID>107</ID>
<type>DE_TO</type>
<position>14.5,-43</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec5</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>13.5,-32</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec6</lparam></gate>
<gate>
<ID>109</ID>
<type>DE_TO</type>
<position>12.5,-43</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec7</lparam></gate>
<gate>
<ID>110</ID>
<type>DA_FROM</type>
<position>59.5,41.5</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec0</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_AND2</type>
<position>-19.5,43.5</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>99 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>DA_FROM</type>
<position>-24.5,44.5</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>113</ID>
<type>DA_FROM</type>
<position>68,-58</position>
<input>
<ID>IN_0</ID>259 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>114</ID>
<type>DA_FROM</type>
<position>-24.5,42.5</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>115</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>20.5,-73.5</position>
<output>
<ID>A_equal_B</ID>176 </output>
<output>
<ID>A_greater_B</ID>174 </output>
<output>
<ID>A_less_B</ID>175 </output>
<input>
<ID>IN_0</ID>177 </input>
<input>
<ID>IN_1</ID>183 </input>
<input>
<ID>IN_2</ID>178 </input>
<input>
<ID>IN_3</ID>184 </input>
<input>
<ID>IN_B_0</ID>180 </input>
<input>
<ID>IN_B_1</ID>181 </input>
<input>
<ID>IN_B_2</ID>179 </input>
<input>
<ID>IN_B_3</ID>182 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>116</ID>
<type>DE_TO</type>
<position>-14.5,43.5</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND0</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_AND2</type>
<position>-19.5,39.5</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>102 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>DA_FROM</type>
<position>74,-47</position>
<input>
<ID>IN_0</ID>246 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>119</ID>
<type>DA_FROM</type>
<position>69,45</position>
<input>
<ID>IN_0</ID>173 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR0</lparam></gate>
<gate>
<ID>120</ID>
<type>DA_FROM</type>
<position>-24.5,40.5</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>121</ID>
<type>DA_FROM</type>
<position>68,-64</position>
<input>
<ID>IN_0</ID>255 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND3</lparam></gate>
<gate>
<ID>122</ID>
<type>DA_FROM</type>
<position>-24.5,38.5</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>123</ID>
<type>DE_TO</type>
<position>-14.5,39.5</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND1</lparam></gate>
<gate>
<ID>124</ID>
<type>DA_FROM</type>
<position>111.5,-28.5</position>
<input>
<ID>IN_0</ID>315 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND6</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_AND2</type>
<position>-19.5,35.5</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>102,-32.5</position>
<input>
<ID>IN_0</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum6</lparam></gate>
<gate>
<ID>127</ID>
<type>DA_FROM</type>
<position>-24.5,36.5</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>128</ID>
<type>DA_FROM</type>
<position>6,-62.5</position>
<input>
<ID>IN_0</ID>187 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>129</ID>
<type>DA_FROM</type>
<position>-24.5,34.5</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>130</ID>
<type>DE_TO</type>
<position>-14.5,35.5</position>
<input>
<ID>IN_0</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND2</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>111.5,-58</position>
<input>
<ID>IN_0</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>7,-67.5</position>
<input>
<ID>IN_0</ID>185 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_AND2</type>
<position>-19.5,31.5</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>DA_FROM</type>
<position>116.5,60</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>-24.5,32.5</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>136</ID>
<type>DA_FROM</type>
<position>0,-67.5</position>
<input>
<ID>IN_0</ID>189 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>137</ID>
<type>DA_FROM</type>
<position>-24.5,30.5</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>138</ID>
<type>DE_TO</type>
<position>-14.5,31.5</position>
<input>
<ID>IN_0</ID>110 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND3</lparam></gate>
<gate>
<ID>139</ID>
<type>DA_FROM</type>
<position>119.5,55</position>
<input>
<ID>IN_0</ID>267 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>140</ID>
<type>DA_FROM</type>
<position>17.5,-62.5</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_AND2</type>
<position>-19.5,27.5</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>DA_FROM</type>
<position>103,39</position>
<input>
<ID>IN_0</ID>272 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum4</lparam></gate>
<gate>
<ID>143</ID>
<type>DA_FROM</type>
<position>-24.5,28.5</position>
<input>
<ID>IN_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>144</ID>
<type>DA_FROM</type>
<position>16.5,-67.5</position>
<input>
<ID>IN_0</ID>178 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>145</ID>
<type>DA_FROM</type>
<position>-24.5,26.5</position>
<input>
<ID>IN_0</ID>111 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>146</ID>
<type>DE_TO</type>
<position>-14.5,27.5</position>
<input>
<ID>IN_0</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND4</lparam></gate>
<gate>
<ID>147</ID>
<type>DA_FROM</type>
<position>111.5,-62</position>
<input>
<ID>IN_0</ID>337 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR7</lparam></gate>
<gate>
<ID>148</ID>
<type>DA_FROM</type>
<position>-24.5,-11.5</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_AND2</type>
<position>-19.5,23.5</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>114 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>DA_FROM</type>
<position>117.5,-47</position>
<input>
<ID>IN_0</ID>326 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>151</ID>
<type>DA_FROM</type>
<position>-24.5,24.5</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>152</ID>
<type>DA_FROM</type>
<position>4,-62.5</position>
<input>
<ID>IN_0</ID>188 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>153</ID>
<type>DA_FROM</type>
<position>-24.5,22.5</position>
<input>
<ID>IN_0</ID>114 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>154</ID>
<type>DE_TO</type>
<position>-14.5,23.5</position>
<input>
<ID>IN_0</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND5</lparam></gate>
<gate>
<ID>155</ID>
<type>AE_SMALL_INVERTER</type>
<position>111.5,38</position>
<input>
<ID>IN_0</ID>271 </input>
<output>
<ID>OUT_0</ID>270 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>156</ID>
<type>DA_FROM</type>
<position>25.5,-67.5</position>
<input>
<ID>IN_0</ID>180 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_AND2</type>
<position>-19.5,19.5</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>158</ID>
<type>DE_TO</type>
<position>122.5,-64.5</position>
<input>
<ID>IN_0</ID>323 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R7</lparam></gate>
<gate>
<ID>159</ID>
<type>DA_FROM</type>
<position>-24.5,20.5</position>
<input>
<ID>IN_0</ID>118 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>160</ID>
<type>DA_FROM</type>
<position>-24.5,18.5</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>161</ID>
<type>DE_TO</type>
<position>-14.5,19.5</position>
<input>
<ID>IN_0</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND6</lparam></gate>
<gate>
<ID>162</ID>
<type>AM_MUX_16x1</type>
<position>118,8</position>
<input>
<ID>IN_0</ID>288 </input>
<input>
<ID>IN_1</ID>288 </input>
<input>
<ID>IN_10</ID>297 </input>
<input>
<ID>IN_11</ID>302 </input>
<input>
<ID>IN_12</ID>300 </input>
<input>
<ID>IN_13</ID>301 </input>
<input>
<ID>IN_14</ID>299 </input>
<input>
<ID>IN_15</ID>298 </input>
<input>
<ID>IN_2</ID>289 </input>
<input>
<ID>IN_3</ID>290 </input>
<input>
<ID>IN_4</ID>292 </input>
<input>
<ID>IN_5</ID>293 </input>
<input>
<ID>IN_6</ID>294 </input>
<input>
<ID>IN_7</ID>294 </input>
<input>
<ID>IN_8</ID>295 </input>
<input>
<ID>IN_9</ID>296 </input>
<output>
<ID>OUT</ID>283 </output>
<input>
<ID>SEL_0</ID>287 </input>
<input>
<ID>SEL_1</ID>286 </input>
<input>
<ID>SEL_2</ID>284 </input>
<input>
<ID>SEL_3</ID>285 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>163</ID>
<type>DA_FROM</type>
<position>-24.5,-19.5</position>
<input>
<ID>IN_0</ID>137 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>164</ID>
<type>AA_AND2</type>
<position>-19.5,15.5</position>
<input>
<ID>IN_0</ID>121 </input>
<input>
<ID>IN_1</ID>120 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_FROM</type>
<position>112.5,47</position>
<input>
<ID>IN_0</ID>280 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>166</ID>
<type>DA_FROM</type>
<position>-24.5,16.5</position>
<input>
<ID>IN_0</ID>121 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>167</ID>
<type>DA_FROM</type>
<position>-24.5,14.5</position>
<input>
<ID>IN_0</ID>120 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>168</ID>
<type>DE_TO</type>
<position>-14.5,15.5</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND7</lparam></gate>
<gate>
<ID>169</ID>
<type>DA_FROM</type>
<position>100.5,-23.5</position>
<input>
<ID>IN_0</ID>321 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>170</ID>
<type>DA_FROM</type>
<position>-24.5,-7.5</position>
<input>
<ID>IN_0</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>171</ID>
<type>DA_FROM</type>
<position>101.5,46</position>
<input>
<ID>IN_0</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>172</ID>
<type>DA_FROM</type>
<position>-24.5,8.5</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>173</ID>
<type>DA_FROM</type>
<position>-24.5,6.5</position>
<input>
<ID>IN_0</ID>123 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>174</ID>
<type>DA_FROM</type>
<position>92,19.5</position>
<input>
<ID>IN_0</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>175</ID>
<type>DA_FROM</type>
<position>-24.5,4.5</position>
<input>
<ID>IN_0</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>176</ID>
<type>DA_FROM</type>
<position>-24.5,2.5</position>
<input>
<ID>IN_0</ID>126 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>177</ID>
<type>DA_FROM</type>
<position>101.5,50</position>
<input>
<ID>IN_0</ID>278 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>178</ID>
<type>DA_FROM</type>
<position>-24.5,-15.5</position>
<input>
<ID>IN_0</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>179</ID>
<type>DA_FROM</type>
<position>-24.5,0.5</position>
<input>
<ID>IN_0</ID>128 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>180</ID>
<type>AE_OR2</type>
<position>-19.5,-0.5</position>
<input>
<ID>IN_0</ID>128 </input>
<input>
<ID>IN_1</ID>127 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>181</ID>
<type>DA_FROM</type>
<position>-24.5,-1.5</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>182</ID>
<type>DA_FROM</type>
<position>-24.5,-3.5</position>
<input>
<ID>IN_0</ID>129 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>183</ID>
<type>AE_OR2</type>
<position>-19.5,-16.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>136 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>184</ID>
<type>DA_FROM</type>
<position>-24.5,-5.5</position>
<input>
<ID>IN_0</ID>130 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>185</ID>
<type>DA_FROM</type>
<position>100.5,-25.5</position>
<input>
<ID>IN_0</ID>322 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>186</ID>
<type>DA_FROM</type>
<position>-24.5,-9.5</position>
<input>
<ID>IN_0</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>187</ID>
<type>AM_MUX_16x1</type>
<position>117,-29</position>
<input>
<ID>IN_0</ID>308 </input>
<input>
<ID>IN_1</ID>308 </input>
<input>
<ID>IN_10</ID>317 </input>
<input>
<ID>IN_11</ID>322 </input>
<input>
<ID>IN_12</ID>320 </input>
<input>
<ID>IN_13</ID>321 </input>
<input>
<ID>IN_14</ID>319 </input>
<input>
<ID>IN_15</ID>318 </input>
<input>
<ID>IN_2</ID>309 </input>
<input>
<ID>IN_3</ID>310 </input>
<input>
<ID>IN_4</ID>312 </input>
<input>
<ID>IN_5</ID>313 </input>
<input>
<ID>IN_6</ID>314 </input>
<input>
<ID>IN_7</ID>314 </input>
<input>
<ID>IN_8</ID>315 </input>
<input>
<ID>IN_9</ID>316 </input>
<output>
<ID>OUT</ID>303 </output>
<input>
<ID>SEL_0</ID>307 </input>
<input>
<ID>SEL_1</ID>306 </input>
<input>
<ID>SEL_2</ID>304 </input>
<input>
<ID>SEL_3</ID>305 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>188</ID>
<type>DA_FROM</type>
<position>-24.5,-13.5</position>
<input>
<ID>IN_0</ID>133 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>189</ID>
<type>DA_FROM</type>
<position>115.5,-47</position>
<input>
<ID>IN_0</ID>325 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>190</ID>
<type>DA_FROM</type>
<position>-24.5,-17.5</position>
<input>
<ID>IN_0</ID>136 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>191</ID>
<type>DA_FROM</type>
<position>91.5,-31.5</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff6</lparam></gate>
<gate>
<ID>192</ID>
<type>DA_FROM</type>
<position>-24.5,-21.5</position>
<input>
<ID>IN_0</ID>138 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>193</ID>
<type>AE_OR2</type>
<position>-19.5,7.5</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>123 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>194</ID>
<type>DA_FROM</type>
<position>111.5,-22.5</position>
<input>
<ID>IN_0</ID>319 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>195</ID>
<type>AE_OR2</type>
<position>-19.5,3.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>140 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>196</ID>
<type>AE_OR2</type>
<position>-19.5,-4.5</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>142 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>197</ID>
<type>AE_OR2</type>
<position>-19.5,-8.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>198</ID>
<type>DA_FROM</type>
<position>118.5,-52</position>
<input>
<ID>IN_0</ID>327 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>199</ID>
<type>AE_OR2</type>
<position>-19.5,-12.5</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>144 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>AE_OR2</type>
<position>-19.5,-20.5</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>DA_FROM</type>
<position>102,-68</position>
<input>
<ID>IN_0</ID>332 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum7</lparam></gate>
<gate>
<ID>202</ID>
<type>DE_TO</type>
<position>-14.5,7.5</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR0</lparam></gate>
<gate>
<ID>203</ID>
<type>DE_TO</type>
<position>-14.5,3.5</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR1</lparam></gate>
<gate>
<ID>204</ID>
<type>DE_TO</type>
<position>-14.5,-0.5</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR2</lparam></gate>
<gate>
<ID>205</ID>
<type>DE_TO</type>
<position>-14.5,-4.5</position>
<input>
<ID>IN_0</ID>142 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR3</lparam></gate>
<gate>
<ID>206</ID>
<type>DA_FROM</type>
<position>100.5,-61</position>
<input>
<ID>IN_0</ID>342 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>207</ID>
<type>DE_TO</type>
<position>-14.5,-8.5</position>
<input>
<ID>IN_0</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR4</lparam></gate>
<gate>
<ID>208</ID>
<type>DE_TO</type>
<position>-14.5,-16.5</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR6</lparam></gate>
<gate>
<ID>209</ID>
<type>DE_TO</type>
<position>-14.5,-20.5</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR7</lparam></gate>
<gate>
<ID>210</ID>
<type>DA_FROM</type>
<position>-24.5,-45.5</position>
<input>
<ID>IN_0</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>211</ID>
<type>DA_FROM</type>
<position>-24.5,-53.5</position>
<input>
<ID>IN_0</ID>160 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>212</ID>
<type>DA_FROM</type>
<position>-24.5,-41.5</position>
<input>
<ID>IN_0</ID>154 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>213</ID>
<type>DA_FROM</type>
<position>-24.5,-25.5</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>214</ID>
<type>DA_FROM</type>
<position>-24.5,-27.5</position>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>215</ID>
<type>DA_FROM</type>
<position>-24.5,-31.5</position>
<input>
<ID>IN_0</ID>162 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>216</ID>
<type>DA_FROM</type>
<position>-24.5,-33.5</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>217</ID>
<type>DA_FROM</type>
<position>-24.5,-37.5</position>
<input>
<ID>IN_0</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>218</ID>
<type>DA_FROM</type>
<position>-24.5,-43.5</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>219</ID>
<type>DA_FROM</type>
<position>-24.5,-51.5</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>220</ID>
<type>DA_FROM</type>
<position>-24.5,-55.5</position>
<input>
<ID>IN_0</ID>159 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>221</ID>
<type>AI_XOR2</type>
<position>-19.5,-26.5</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>148 </input>
<output>
<ID>OUT</ID>163 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>AI_XOR2</type>
<position>-19.5,-30.5</position>
<input>
<ID>IN_0</ID>161 </input>
<input>
<ID>IN_1</ID>162 </input>
<output>
<ID>OUT</ID>164 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>223</ID>
<type>AI_XOR2</type>
<position>-19.5,-34.5</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>149 </input>
<output>
<ID>OUT</ID>165 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>224</ID>
<type>AI_XOR2</type>
<position>-19.5,-38.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>152 </input>
<output>
<ID>OUT</ID>166 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>225</ID>
<type>AI_XOR2</type>
<position>-19.5,-42.5</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>153 </input>
<output>
<ID>OUT</ID>167 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>226</ID>
<type>AI_XOR2</type>
<position>-19.5,-46.5</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>155 </input>
<output>
<ID>OUT</ID>168 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>AI_XOR2</type>
<position>-19.5,-50.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>157 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>AI_XOR2</type>
<position>-19.5,-54.5</position>
<input>
<ID>IN_0</ID>160 </input>
<input>
<ID>IN_1</ID>159 </input>
<output>
<ID>OUT</ID>170 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>229</ID>
<type>DE_TO</type>
<position>-14.5,-26.5</position>
<input>
<ID>IN_0</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR0</lparam></gate>
<gate>
<ID>230</ID>
<type>DE_TO</type>
<position>-14.5,-30.5</position>
<input>
<ID>IN_0</ID>164 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR1</lparam></gate>
<gate>
<ID>231</ID>
<type>DE_TO</type>
<position>-14.5,-34.5</position>
<input>
<ID>IN_0</ID>165 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR2</lparam></gate>
<gate>
<ID>232</ID>
<type>DE_TO</type>
<position>-14.5,-38.5</position>
<input>
<ID>IN_0</ID>166 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR3</lparam></gate>
<gate>
<ID>233</ID>
<type>DE_TO</type>
<position>-14.5,-42.5</position>
<input>
<ID>IN_0</ID>167 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR4</lparam></gate>
<gate>
<ID>234</ID>
<type>DA_FROM</type>
<position>57,-23.5</position>
<input>
<ID>IN_0</ID>241 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>235</ID>
<type>DE_TO</type>
<position>-14.5,-46.5</position>
<input>
<ID>IN_0</ID>168 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR5</lparam></gate>
<gate>
<ID>236</ID>
<type>DE_TO</type>
<position>-14.5,-50.5</position>
<input>
<ID>IN_0</ID>169 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR6</lparam></gate>
<gate>
<ID>237</ID>
<type>DE_TO</type>
<position>-14.5,-54.5</position>
<input>
<ID>IN_0</ID>170 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR7</lparam></gate>
<gate>
<ID>238</ID>
<type>DE_TO</type>
<position>79,-64.5</position>
<input>
<ID>IN_0</ID>243 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R3</lparam></gate>
<gate>
<ID>239</ID>
<type>DA_FROM</type>
<position>69,43</position>
<input>
<ID>IN_0</ID>171 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND0</lparam></gate>
<gate>
<ID>240</ID>
<type>DA_FROM</type>
<position>58,44</position>
<input>
<ID>IN_0</ID>172 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR0</lparam></gate>
<gate>
<ID>241</ID>
<type>DA_FROM</type>
<position>68,-62</position>
<input>
<ID>IN_0</ID>257 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR3</lparam></gate>
<gate>
<ID>242</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>2,-73.5</position>
<output>
<ID>A_equal_B</ID>194 </output>
<output>
<ID>A_greater_B</ID>195 </output>
<output>
<ID>A_less_B</ID>193 </output>
<input>
<ID>IN_0</ID>189 </input>
<input>
<ID>IN_1</ID>192 </input>
<input>
<ID>IN_2</ID>190 </input>
<input>
<ID>IN_3</ID>191 </input>
<input>
<ID>IN_B_0</ID>185 </input>
<input>
<ID>IN_B_1</ID>187 </input>
<input>
<ID>IN_B_2</ID>186 </input>
<input>
<ID>IN_B_3</ID>188 </input>
<input>
<ID>in_A_equal_B</ID>176 </input>
<input>
<ID>in_A_greater_B</ID>174 </input>
<input>
<ID>in_A_less_B</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>243</ID>
<type>DA_FROM</type>
<position>22.5,-62.5</position>
<input>
<ID>IN_0</ID>182 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>244</ID>
<type>DA_FROM</type>
<position>118.5,25.5</position>
<input>
<ID>IN_0</ID>286 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>245</ID>
<type>DA_FROM</type>
<position>23.5,-67.5</position>
<input>
<ID>IN_0</ID>179 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>246</ID>
<type>DA_FROM</type>
<position>-2,-67.5</position>
<input>
<ID>IN_0</ID>190 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>247</ID>
<type>DA_FROM</type>
<position>118.5,-16.5</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>248</ID>
<type>DA_FROM</type>
<position>-1,-62.5</position>
<input>
<ID>IN_0</ID>192 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>249</ID>
<type>AE_SMALL_INVERTER</type>
<position>107,2.5</position>
<input>
<ID>IN_0</ID>288 </input>
<output>
<ID>OUT_0</ID>289 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>250</ID>
<type>DA_FROM</type>
<position>-3,-62.5</position>
<input>
<ID>IN_0</ID>191 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>251</ID>
<type>DA_FROM</type>
<position>18.5,-67.5</position>
<input>
<ID>IN_0</ID>177 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>252</ID>
<type>DA_FROM</type>
<position>103,7</position>
<input>
<ID>IN_0</ID>294 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec5</lparam></gate>
<gate>
<ID>253</ID>
<type>DA_FROM</type>
<position>24.5,-62.5</position>
<input>
<ID>IN_0</ID>181 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>254</ID>
<type>DA_FROM</type>
<position>15.5,-62.5</position>
<input>
<ID>IN_0</ID>184 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>255</ID>
<type>DA_FROM</type>
<position>91.5,-67</position>
<input>
<ID>IN_0</ID>333 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff7</lparam></gate>
<gate>
<ID>256</ID>
<type>DA_FROM</type>
<position>5,-67.5</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>257</ID>
<type>DE_TO</type>
<position>-8,-71.5</position>
<input>
<ID>IN_0</ID>195 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>258</ID>
<type>DA_FROM</type>
<position>102,-30</position>
<input>
<ID>IN_0</ID>314 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec6</lparam></gate>
<gate>
<ID>259</ID>
<type>DE_TO</type>
<position>-11,-73.5</position>
<input>
<ID>IN_0</ID>194 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>260</ID>
<type>DE_TO</type>
<position>-8,-75.5</position>
<input>
<ID>IN_0</ID>193 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>261</ID>
<type>DA_FROM</type>
<position>116.5,-16.5</position>
<input>
<ID>IN_0</ID>304 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>262</ID>
<type>AE_OR2</type>
<position>-19,-71.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>195 </input>
<output>
<ID>OUT</ID>196 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>263</ID>
<type>AE_OR2</type>
<position>-19,-75.5</position>
<input>
<ID>IN_0</ID>193 </input>
<input>
<ID>IN_1</ID>194 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>264</ID>
<type>DA_FROM</type>
<position>112.5,45</position>
<input>
<ID>IN_0</ID>277 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR4</lparam></gate>
<gate>
<ID>265</ID>
<type>DE_TO</type>
<position>-24,-71.5</position>
<input>
<ID>IN_0</ID>196 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>266</ID>
<type>DE_TO</type>
<position>-24,-75.5</position>
<input>
<ID>IN_0</ID>197 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>267</ID>
<type>DA_FROM</type>
<position>118.5,60</position>
<input>
<ID>IN_0</ID>266 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>268</ID>
<type>DA_FROM</type>
<position>69,47</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>269</ID>
<type>DA_FROM</type>
<position>117.5,20.5</position>
<input>
<ID>IN_0</ID>284 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>270</ID>
<type>DA_FROM</type>
<position>69,49</position>
<input>
<ID>IN_0</ID>199 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>271</ID>
<type>DA_FROM</type>
<position>112.5,49</position>
<input>
<ID>IN_0</ID>279 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>272</ID>
<type>DA_FROM</type>
<position>58,48</position>
<input>
<ID>IN_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>273</ID>
<type>AE_SMALL_INVERTER</type>
<position>111.5,3.5</position>
<input>
<ID>IN_0</ID>291 </input>
<output>
<ID>OUT_0</ID>290 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>274</ID>
<type>DA_FROM</type>
<position>58,50</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>275</ID>
<type>DA_FROM</type>
<position>92.5,40</position>
<input>
<ID>IN_0</ID>273 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff4</lparam></gate>
<gate>
<ID>276</ID>
<type>DA_FROM</type>
<position>58,46</position>
<input>
<ID>IN_0</ID>202 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>277</ID>
<type>DA_FROM</type>
<position>48.5,21.5</position>
<input>
<ID>IN_0</ID>208 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>278</ID>
<type>DE_TO</type>
<position>80,8</position>
<input>
<ID>IN_0</ID>203 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1</lparam></gate>
<gate>
<ID>279</ID>
<type>AM_MUX_16x1</type>
<position>74.5,8</position>
<input>
<ID>IN_0</ID>208 </input>
<input>
<ID>IN_1</ID>208 </input>
<input>
<ID>IN_10</ID>217 </input>
<input>
<ID>IN_11</ID>222 </input>
<input>
<ID>IN_12</ID>220 </input>
<input>
<ID>IN_13</ID>221 </input>
<input>
<ID>IN_14</ID>219 </input>
<input>
<ID>IN_15</ID>218 </input>
<input>
<ID>IN_2</ID>209 </input>
<input>
<ID>IN_3</ID>210 </input>
<input>
<ID>IN_4</ID>212 </input>
<input>
<ID>IN_5</ID>213 </input>
<input>
<ID>IN_6</ID>214 </input>
<input>
<ID>IN_7</ID>214 </input>
<input>
<ID>IN_8</ID>215 </input>
<input>
<ID>IN_9</ID>216 </input>
<output>
<ID>OUT</ID>203 </output>
<input>
<ID>SEL_0</ID>207 </input>
<input>
<ID>SEL_1</ID>206 </input>
<input>
<ID>SEL_2</ID>204 </input>
<input>
<ID>SEL_3</ID>205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>280</ID>
<type>DA_FROM</type>
<position>48.5,19.5</position>
<input>
<ID>IN_0</ID>211 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>281</ID>
<type>DA_FROM</type>
<position>76,20.5</position>
<input>
<ID>IN_0</ID>207 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>282</ID>
<type>DA_FROM</type>
<position>75,25.5</position>
<input>
<ID>IN_0</ID>206 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>283</ID>
<type>DA_FROM</type>
<position>74,20.5</position>
<input>
<ID>IN_0</ID>204 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>284</ID>
<type>DA_FROM</type>
<position>73,25.5</position>
<input>
<ID>IN_0</ID>205 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>285</ID>
<type>DA_FROM</type>
<position>47.5,-53</position>
<input>
<ID>IN_0</ID>251 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>286</ID>
<type>AE_SMALL_INVERTER</type>
<position>63.5,2.5</position>
<input>
<ID>IN_0</ID>208 </input>
<output>
<ID>OUT_0</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>287</ID>
<type>AE_SMALL_INVERTER</type>
<position>68,3.5</position>
<input>
<ID>IN_0</ID>211 </input>
<output>
<ID>OUT_0</ID>210 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>288</ID>
<type>DA_FROM</type>
<position>59.5,4.5</position>
<input>
<ID>IN_0</ID>212 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum1</lparam></gate>
<gate>
<ID>289</ID>
<type>DA_FROM</type>
<position>49,5.5</position>
<input>
<ID>IN_0</ID>213 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff1</lparam></gate>
<gate>
<ID>290</ID>
<type>DA_FROM</type>
<position>59.5,7</position>
<input>
<ID>IN_0</ID>214 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec1</lparam></gate>
<gate>
<ID>291</ID>
<type>DA_FROM</type>
<position>69,10.5</position>
<input>
<ID>IN_0</ID>217 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR1</lparam></gate>
<gate>
<ID>292</ID>
<type>DA_FROM</type>
<position>69,8.5</position>
<input>
<ID>IN_0</ID>215 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND1</lparam></gate>
<gate>
<ID>293</ID>
<type>DA_FROM</type>
<position>58,9.5</position>
<input>
<ID>IN_0</ID>216 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR1</lparam></gate>
<gate>
<ID>294</ID>
<type>DA_FROM</type>
<position>48,-67</position>
<input>
<ID>IN_0</ID>253 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff3</lparam></gate>
<gate>
<ID>295</ID>
<type>DA_FROM</type>
<position>69,12.5</position>
<input>
<ID>IN_0</ID>220 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>296</ID>
<type>DA_FROM</type>
<position>69,14.5</position>
<input>
<ID>IN_0</ID>219 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>297</ID>
<type>DA_FROM</type>
<position>58,13.5</position>
<input>
<ID>IN_0</ID>221 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>298</ID>
<type>DA_FROM</type>
<position>57,-25.5</position>
<input>
<ID>IN_0</ID>242 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>299</ID>
<type>DA_FROM</type>
<position>58,11.5</position>
<input>
<ID>IN_0</ID>222 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>300</ID>
<type>DA_FROM</type>
<position>47.5,-15.5</position>
<input>
<ID>IN_0</ID>228 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>301</ID>
<type>DE_TO</type>
<position>79,-29</position>
<input>
<ID>IN_0</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R2</lparam></gate>
<gate>
<ID>302</ID>
<type>AM_MUX_16x1</type>
<position>73.5,-29</position>
<input>
<ID>IN_0</ID>228 </input>
<input>
<ID>IN_1</ID>228 </input>
<input>
<ID>IN_10</ID>237 </input>
<input>
<ID>IN_11</ID>242 </input>
<input>
<ID>IN_12</ID>240 </input>
<input>
<ID>IN_13</ID>241 </input>
<input>
<ID>IN_14</ID>239 </input>
<input>
<ID>IN_15</ID>238 </input>
<input>
<ID>IN_2</ID>229 </input>
<input>
<ID>IN_3</ID>230 </input>
<input>
<ID>IN_4</ID>232 </input>
<input>
<ID>IN_5</ID>233 </input>
<input>
<ID>IN_6</ID>234 </input>
<input>
<ID>IN_7</ID>234 </input>
<input>
<ID>IN_8</ID>235 </input>
<input>
<ID>IN_9</ID>236 </input>
<output>
<ID>OUT</ID>223 </output>
<input>
<ID>SEL_0</ID>227 </input>
<input>
<ID>SEL_1</ID>226 </input>
<input>
<ID>SEL_2</ID>224 </input>
<input>
<ID>SEL_3</ID>225 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>303</ID>
<type>DA_FROM</type>
<position>57,-57</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>304</ID>
<type>DA_FROM</type>
<position>47.5,-17.5</position>
<input>
<ID>IN_0</ID>231 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>305</ID>
<type>DA_FROM</type>
<position>74,-11.5</position>
<input>
<ID>IN_0</ID>226 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>306</ID>
<type>DA_FROM</type>
<position>72,-47</position>
<input>
<ID>IN_0</ID>245 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>307</ID>
<type>DA_FROM</type>
<position>72,-11.5</position>
<input>
<ID>IN_0</ID>225 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>308</ID>
<type>AE_SMALL_INVERTER</type>
<position>62.5,-34.5</position>
<input>
<ID>IN_0</ID>228 </input>
<output>
<ID>OUT_0</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>309</ID>
<type>AE_SMALL_INVERTER</type>
<position>67,-33.5</position>
<input>
<ID>IN_0</ID>231 </input>
<output>
<ID>OUT_0</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>310</ID>
<type>DA_FROM</type>
<position>92,54</position>
<input>
<ID>IN_0</ID>271 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>311</ID>
<type>DA_FROM</type>
<position>48,-31.5</position>
<input>
<ID>IN_0</ID>233 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff2</lparam></gate>
<gate>
<ID>312</ID>
<type>DA_FROM</type>
<position>68,-26.5</position>
<input>
<ID>IN_0</ID>237 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR2</lparam></gate>
<gate>
<ID>313</ID>
<type>DA_FROM</type>
<position>57,-63</position>
<input>
<ID>IN_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR3</lparam></gate>
<gate>
<ID>314</ID>
<type>DA_FROM</type>
<position>57,-27.5</position>
<input>
<ID>IN_0</ID>236 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR2</lparam></gate>
<gate>
<ID>315</ID>
<type>DA_FROM</type>
<position>68,-22.5</position>
<input>
<ID>IN_0</ID>239 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>316</ID>
<type>DA_FROM</type>
<position>57,-21.5</position>
<input>
<ID>IN_0</ID>238 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>317</ID>
<type>DA_FROM</type>
<position>47.5,-51</position>
<input>
<ID>IN_0</ID>248 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>318</ID>
<type>AM_MUX_16x1</type>
<position>73.5,-64.5</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>248 </input>
<input>
<ID>IN_10</ID>257 </input>
<input>
<ID>IN_11</ID>262 </input>
<input>
<ID>IN_12</ID>260 </input>
<input>
<ID>IN_13</ID>261 </input>
<input>
<ID>IN_14</ID>259 </input>
<input>
<ID>IN_15</ID>258 </input>
<input>
<ID>IN_2</ID>249 </input>
<input>
<ID>IN_3</ID>250 </input>
<input>
<ID>IN_4</ID>252 </input>
<input>
<ID>IN_5</ID>253 </input>
<input>
<ID>IN_6</ID>254 </input>
<input>
<ID>IN_7</ID>254 </input>
<input>
<ID>IN_8</ID>255 </input>
<input>
<ID>IN_9</ID>256 </input>
<output>
<ID>OUT</ID>243 </output>
<input>
<ID>SEL_0</ID>247 </input>
<input>
<ID>SEL_1</ID>246 </input>
<input>
<ID>SEL_2</ID>244 </input>
<input>
<ID>SEL_3</ID>245 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>319</ID>
<type>DA_FROM</type>
<position>75,-52</position>
<input>
<ID>IN_0</ID>247 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>320</ID>
<type>DA_FROM</type>
<position>73,-52</position>
<input>
<ID>IN_0</ID>244 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>321</ID>
<type>AE_SMALL_INVERTER</type>
<position>62.5,-70</position>
<input>
<ID>IN_0</ID>248 </input>
<output>
<ID>OUT_0</ID>249 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>322</ID>
<type>AE_SMALL_INVERTER</type>
<position>67,-69</position>
<input>
<ID>IN_0</ID>251 </input>
<output>
<ID>OUT_0</ID>250 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>323</ID>
<type>DA_FROM</type>
<position>58.5,-68</position>
<input>
<ID>IN_0</ID>252 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum3</lparam></gate>
<gate>
<ID>324</ID>
<type>DA_FROM</type>
<position>58.5,-65.5</position>
<input>
<ID>IN_0</ID>254 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec3</lparam></gate>
<gate>
<ID>325</ID>
<type>DA_FROM</type>
<position>68,-60</position>
<input>
<ID>IN_0</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>326</ID>
<type>DA_FROM</type>
<position>57,-59</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>327</ID>
<type>DA_FROM</type>
<position>57,-61</position>
<input>
<ID>IN_0</ID>262 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>328</ID>
<type>DA_FROM</type>
<position>92,56</position>
<input>
<ID>IN_0</ID>268 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>329</ID>
<type>DE_TO</type>
<position>123.5,42.5</position>
<input>
<ID>IN_0</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R4</lparam></gate>
<gate>
<ID>330</ID>
<type>DA_FROM</type>
<position>101.5,15.5</position>
<input>
<ID>IN_0</ID>298 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>331</ID>
<type>AM_MUX_16x1</type>
<position>118,42.5</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>268 </input>
<input>
<ID>IN_10</ID>277 </input>
<input>
<ID>IN_11</ID>282 </input>
<input>
<ID>IN_12</ID>280 </input>
<input>
<ID>IN_13</ID>281 </input>
<input>
<ID>IN_14</ID>279 </input>
<input>
<ID>IN_15</ID>278 </input>
<input>
<ID>IN_2</ID>269 </input>
<input>
<ID>IN_3</ID>270 </input>
<input>
<ID>IN_4</ID>272 </input>
<input>
<ID>IN_5</ID>273 </input>
<input>
<ID>IN_6</ID>274 </input>
<input>
<ID>IN_7</ID>274 </input>
<input>
<ID>IN_8</ID>275 </input>
<input>
<ID>IN_9</ID>276 </input>
<output>
<ID>OUT</ID>263 </output>
<input>
<ID>SEL_0</ID>267 </input>
<input>
<ID>SEL_1</ID>266 </input>
<input>
<ID>SEL_2</ID>264 </input>
<input>
<ID>SEL_3</ID>265 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>332</ID>
<type>DA_FROM</type>
<position>111.5,-24.5</position>
<input>
<ID>IN_0</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>333</ID>
<type>DA_FROM</type>
<position>117.5,55</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>334</ID>
<type>AE_SMALL_INVERTER</type>
<position>107,37</position>
<input>
<ID>IN_0</ID>268 </input>
<output>
<ID>OUT_0</ID>269 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>335</ID>
<type>DA_FROM</type>
<position>103,41.5</position>
<input>
<ID>IN_0</ID>274 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec4</lparam></gate>
<gate>
<ID>336</ID>
<type>DA_FROM</type>
<position>111.5,-64</position>
<input>
<ID>IN_0</ID>335 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND7</lparam></gate>
<gate>
<ID>337</ID>
<type>DA_FROM</type>
<position>112.5,43</position>
<input>
<ID>IN_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND4</lparam></gate>
<gate>
<ID>338</ID>
<type>DA_FROM</type>
<position>101.5,44</position>
<input>
<ID>IN_0</ID>276 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR4</lparam></gate>
<gate>
<ID>339</ID>
<type>DA_FROM</type>
<position>101.5,48</position>
<input>
<ID>IN_0</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>340</ID>
<type>DA_FROM</type>
<position>92,21.5</position>
<input>
<ID>IN_0</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>341</ID>
<type>DE_TO</type>
<position>123.5,8</position>
<input>
<ID>IN_0</ID>283 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R5</lparam></gate>
<gate>
<ID>342</ID>
<type>DA_FROM</type>
<position>119.5,20.5</position>
<input>
<ID>IN_0</ID>287 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>343</ID>
<type>DA_FROM</type>
<position>116.5,25.5</position>
<input>
<ID>IN_0</ID>285 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>344</ID>
<type>DA_FROM</type>
<position>91,-53</position>
<input>
<ID>IN_0</ID>331 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>345</ID>
<type>DA_FROM</type>
<position>103,4.5</position>
<input>
<ID>IN_0</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum5</lparam></gate>
<gate>
<ID>346</ID>
<type>DA_FROM</type>
<position>92.5,5.5</position>
<input>
<ID>IN_0</ID>293 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff5</lparam></gate>
<gate>
<ID>347</ID>
<type>DA_FROM</type>
<position>112.5,10.5</position>
<input>
<ID>IN_0</ID>297 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR5</lparam></gate>
<gate>
<ID>348</ID>
<type>DA_FROM</type>
<position>112.5,8.5</position>
<input>
<ID>IN_0</ID>295 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND5</lparam></gate>
<gate>
<ID>349</ID>
<type>DA_FROM</type>
<position>101.5,9.5</position>
<input>
<ID>IN_0</ID>296 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR5</lparam></gate>
<gate>
<ID>350</ID>
<type>DA_FROM</type>
<position>112.5,12.5</position>
<input>
<ID>IN_0</ID>300 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>351</ID>
<type>DA_FROM</type>
<position>112.5,14.5</position>
<input>
<ID>IN_0</ID>299 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>352</ID>
<type>DA_FROM</type>
<position>101.5,13.5</position>
<input>
<ID>IN_0</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>353</ID>
<type>DA_FROM</type>
<position>101.5,11.5</position>
<input>
<ID>IN_0</ID>302 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>354</ID>
<type>DA_FROM</type>
<position>91,-15.5</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>355</ID>
<type>DE_TO</type>
<position>122.5,-29</position>
<input>
<ID>IN_0</ID>303 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R6</lparam></gate>
<gate>
<ID>356</ID>
<type>DA_FROM</type>
<position>100.5,-57</position>
<input>
<ID>IN_0</ID>338 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>357</ID>
<type>DA_FROM</type>
<position>91,-17.5</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>358</ID>
<type>DA_FROM</type>
<position>117.5,-11.5</position>
<input>
<ID>IN_0</ID>306 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>359</ID>
<type>DA_FROM</type>
<position>115.5,-11.5</position>
<input>
<ID>IN_0</ID>305 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>360</ID>
<type>AE_SMALL_INVERTER</type>
<position>106,-34.5</position>
<input>
<ID>IN_0</ID>308 </input>
<output>
<ID>OUT_0</ID>309 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>361</ID>
<type>AE_SMALL_INVERTER</type>
<position>110.5,-33.5</position>
<input>
<ID>IN_0</ID>311 </input>
<output>
<ID>OUT_0</ID>310 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>362</ID>
<type>DA_FROM</type>
<position>111.5,-26.5</position>
<input>
<ID>IN_0</ID>317 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR6</lparam></gate>
<gate>
<ID>363</ID>
<type>DA_FROM</type>
<position>100.5,-63</position>
<input>
<ID>IN_0</ID>336 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR7</lparam></gate>
<gate>
<ID>364</ID>
<type>DA_FROM</type>
<position>100.5,-27.5</position>
<input>
<ID>IN_0</ID>316 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR6</lparam></gate>
<gate>
<ID>365</ID>
<type>DA_FROM</type>
<position>100.5,-21.5</position>
<input>
<ID>IN_0</ID>318 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>366</ID>
<type>DA_FROM</type>
<position>91,-51</position>
<input>
<ID>IN_0</ID>328 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>367</ID>
<type>AM_MUX_16x1</type>
<position>117,-64.5</position>
<input>
<ID>IN_0</ID>328 </input>
<input>
<ID>IN_1</ID>328 </input>
<input>
<ID>IN_10</ID>337 </input>
<input>
<ID>IN_11</ID>342 </input>
<input>
<ID>IN_12</ID>340 </input>
<input>
<ID>IN_13</ID>341 </input>
<input>
<ID>IN_14</ID>339 </input>
<input>
<ID>IN_15</ID>338 </input>
<input>
<ID>IN_2</ID>329 </input>
<input>
<ID>IN_3</ID>330 </input>
<input>
<ID>IN_4</ID>332 </input>
<input>
<ID>IN_5</ID>333 </input>
<input>
<ID>IN_6</ID>334 </input>
<input>
<ID>IN_7</ID>334 </input>
<input>
<ID>IN_8</ID>335 </input>
<input>
<ID>IN_9</ID>336 </input>
<output>
<ID>OUT</ID>323 </output>
<input>
<ID>SEL_0</ID>327 </input>
<input>
<ID>SEL_1</ID>326 </input>
<input>
<ID>SEL_2</ID>324 </input>
<input>
<ID>SEL_3</ID>325 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>368</ID>
<type>DA_FROM</type>
<position>116.5,-52</position>
<input>
<ID>IN_0</ID>324 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>369</ID>
<type>AE_SMALL_INVERTER</type>
<position>106,-70</position>
<input>
<ID>IN_0</ID>328 </input>
<output>
<ID>OUT_0</ID>329 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>370</ID>
<type>AE_SMALL_INVERTER</type>
<position>110.5,-69</position>
<input>
<ID>IN_0</ID>331 </input>
<output>
<ID>OUT_0</ID>330 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>371</ID>
<type>DA_FROM</type>
<position>102,-65.5</position>
<input>
<ID>IN_0</ID>334 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec7</lparam></gate>
<gate>
<ID>372</ID>
<type>DA_FROM</type>
<position>111.5,-60</position>
<input>
<ID>IN_0</ID>340 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>373</ID>
<type>DA_FROM</type>
<position>100.5,-59</position>
<input>
<ID>IN_0</ID>341 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>77.5,42.5,78,42.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<connection>
<GID>5</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>74,52,74,53</points>
<connection>
<GID>8</GID>
<name>SEL_2</name></connection>
<connection>
<GID>16</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,52,73,58</points>
<connection>
<GID>8</GID>
<name>SEL_3</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,52,75,58</points>
<connection>
<GID>8</GID>
<name>SEL_1</name></connection>
<connection>
<GID>15</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>76,52,76,53</points>
<connection>
<GID>8</GID>
<name>SEL_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,38.5,23.5,38.5</points>
<connection>
<GID>70</GID>
<name>carry_in</name></connection>
<connection>
<GID>69</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>40,41.5,40,42.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>41.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>36.5,41.5,40,41.5</points>
<connection>
<GID>69</GID>
<name>IN_B_0</name></connection>
<intersection>40 1</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,41.5,35.5,42</points>
<connection>
<GID>69</GID>
<name>IN_B_1</name></connection>
<intersection>42 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>38,42,38,42.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35.5,42,38,42</points>
<intersection>35.5 0</intersection>
<intersection>38 1</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,41.5,34.5,42.5</points>
<connection>
<GID>69</GID>
<name>IN_B_2</name></connection>
<intersection>42.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>34.5,42.5,36,42.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>33.5,41.5,33.5,42.5</points>
<connection>
<GID>69</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>72</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,41.5,29.5,42</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>42 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>31,42,31,42.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>29.5,42,31,42</points>
<intersection>29.5 0</intersection>
<intersection>31 1</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,41.5,28.5,42</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>42 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>29,42,29,42.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,42,29,42</points>
<intersection>28.5 0</intersection>
<intersection>29 1</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,41.5,27.5,42</points>
<connection>
<GID>69</GID>
<name>IN_2</name></connection>
<intersection>42 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>27,42,27,42.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27,42,27.5,42</points>
<intersection>27 1</intersection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,42,25,42.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>42 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>26.5,41.5,26.5,42</points>
<connection>
<GID>69</GID>
<name>IN_3</name></connection>
<intersection>42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>25,42,26.5,42</points>
<intersection>25 0</intersection>
<intersection>26.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>22,41.5,22,42.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>41.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>19,41.5,22,41.5</points>
<connection>
<GID>70</GID>
<name>IN_B_0</name></connection>
<intersection>22 1</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,41.5,18,42</points>
<connection>
<GID>70</GID>
<name>IN_B_1</name></connection>
<intersection>42 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>20,42,20,42.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>18,42,20,42</points>
<intersection>18 0</intersection>
<intersection>20 1</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,41.5,17,42.5</points>
<connection>
<GID>70</GID>
<name>IN_B_2</name></connection>
<intersection>42.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>17,42.5,18,42.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,41.5,16,42.5</points>
<connection>
<GID>70</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>22</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,41.5,12,42</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>42 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>13,42,13,42.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>12,42,13,42</points>
<intersection>12 0</intersection>
<intersection>13 1</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,41.5,11,42.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,42,9,42.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>42 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>10,41.5,10,42</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>9,42,10,42</points>
<intersection>9 0</intersection>
<intersection>10 1</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,41.5,7,42.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>41.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>7,41.5,9,41.5</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,32.5,34.5,33</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>33 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>33,33,33,33.5</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>33,33,34.5,33</points>
<intersection>33 1</intersection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,33,32,33.5</points>
<connection>
<GID>69</GID>
<name>OUT_1</name></connection>
<intersection>33 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>32.5,32.5,32.5,33</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32,33,32.5,33</points>
<intersection>32 0</intersection>
<intersection>32.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,33,31,33.5</points>
<connection>
<GID>69</GID>
<name>OUT_2</name></connection>
<intersection>33 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>30.5,32.5,30.5,33</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30.5,33,31,33</points>
<intersection>30.5 1</intersection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,32.5,28.5,33</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>33 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>30,33,30,33.5</points>
<connection>
<GID>69</GID>
<name>OUT_3</name></connection>
<intersection>33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,33,30,33</points>
<intersection>28.5 0</intersection>
<intersection>30 1</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,33,15.5,33.5</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>33 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>17,32.5,17,33</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>15.5,33,17,33</points>
<intersection>15.5 0</intersection>
<intersection>17 1</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,32.5,15,33</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>33 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>14.5,33,14.5,33.5</points>
<connection>
<GID>70</GID>
<name>OUT_1</name></connection>
<intersection>33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>14.5,33,15,33</points>
<intersection>14.5 1</intersection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,32.5,13,33</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>33 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>13.5,33,13.5,33.5</points>
<connection>
<GID>70</GID>
<name>OUT_2</name></connection>
<intersection>33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>13,33,13.5,33</points>
<intersection>13 0</intersection>
<intersection>13.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,32.5,11,33</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>33 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>12.5,33,12.5,33.5</points>
<connection>
<GID>70</GID>
<name>OUT_3</name></connection>
<intersection>33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11,33,12.5,33</points>
<intersection>11 0</intersection>
<intersection>12.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,38.5,40.5,38.5</points>
<connection>
<GID>69</GID>
<name>carry_in</name></connection>
<intersection>40.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>40.5,38,40.5,38.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>38.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,32,6,36.5</points>
<connection>
<GID>70</GID>
<name>overflow</name></connection>
<intersection>32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>6,32,7.5,32</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,32,5.5,38.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,38.5,6,38.5</points>
<connection>
<GID>70</GID>
<name>carry_out</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,6,23.5,6</points>
<connection>
<GID>53</GID>
<name>carry_in</name></connection>
<connection>
<GID>52</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,9,29.5,9.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>9.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>31,9.5,31,10</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>9.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>29.5,9.5,31,9.5</points>
<intersection>29.5 0</intersection>
<intersection>31 1</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,9,28.5,9.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>9.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>29,9.5,29,10</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>9.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,9.5,29,9.5</points>
<intersection>28.5 0</intersection>
<intersection>29 1</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,9,27.5,9.5</points>
<connection>
<GID>52</GID>
<name>IN_2</name></connection>
<intersection>9.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>27,9.5,27,10</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>9.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27,9.5,27.5,9.5</points>
<intersection>27 1</intersection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,9.5,25,10</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>9.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>26.5,9,26.5,9.5</points>
<connection>
<GID>52</GID>
<name>IN_3</name></connection>
<intersection>9.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>25,9.5,26.5,9.5</points>
<intersection>25 0</intersection>
<intersection>26.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,9,12,9.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>9.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>13,9.5,13,10</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>9.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>12,9.5,13,9.5</points>
<intersection>12 0</intersection>
<intersection>13 1</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,9,11,10</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,9.5,9,10</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>9.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>10,9,10,9.5</points>
<connection>
<GID>53</GID>
<name>IN_2</name></connection>
<intersection>9.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>9,9.5,10,9.5</points>
<intersection>9 0</intersection>
<intersection>10 1</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,9,7,10</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>9 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>7,9,9,9</points>
<connection>
<GID>53</GID>
<name>IN_3</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,0,34.5,0.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>33,0.5,33,1</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>33,0.5,34.5,0.5</points>
<intersection>33 1</intersection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,0.5,32,1</points>
<connection>
<GID>52</GID>
<name>OUT_1</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>32.5,0,32.5,0.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32,0.5,32.5,0.5</points>
<intersection>32 0</intersection>
<intersection>32.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,0.5,31,1</points>
<connection>
<GID>52</GID>
<name>OUT_2</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>30.5,0,30.5,0.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30.5,0.5,31,0.5</points>
<intersection>30.5 1</intersection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,0,28.5,0.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>30,0.5,30,1</points>
<connection>
<GID>52</GID>
<name>OUT_3</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,0.5,30,0.5</points>
<intersection>28.5 0</intersection>
<intersection>30 1</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,0.5,15.5,1</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>17,0,17,0.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>15.5,0.5,17,0.5</points>
<intersection>15.5 0</intersection>
<intersection>17 1</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,0,15,0.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>14.5,0.5,14.5,1</points>
<connection>
<GID>53</GID>
<name>OUT_1</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>14.5,0.5,15,0.5</points>
<intersection>14.5 1</intersection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,0,13,0.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>13.5,0.5,13.5,1</points>
<connection>
<GID>53</GID>
<name>OUT_2</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>13,0.5,13.5,0.5</points>
<intersection>13 0</intersection>
<intersection>13.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,0,11,0.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>12.5,0.5,12.5,1</points>
<connection>
<GID>53</GID>
<name>OUT_3</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11,0.5,12.5,0.5</points>
<intersection>11 0</intersection>
<intersection>12.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-0.5,6,4</points>
<connection>
<GID>53</GID>
<name>overflow</name></connection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>6,-0.5,7.5,-0.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-0.5,5.5,6</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,6,6,6</points>
<connection>
<GID>53</GID>
<name>carry_out</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>33.5,9,33.5,9.5</points>
<connection>
<GID>52</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>35.5,9,35.5,9.5</points>
<connection>
<GID>52</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>62</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>34.5,9,34.5,9.5</points>
<connection>
<GID>52</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>62</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>36.5,9,36.5,9.5</points>
<connection>
<GID>52</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>62</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,13.5,33.5,15</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,13.5,34.5,15</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>15 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>34.5,15,35.5,15</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>36.5,13.5,39.5,13.5</points>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<intersection>39.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>39.5,13.5,39.5,15</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>13.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,13.5,35.5,14</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<intersection>14 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>37.5,14,37.5,15</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35.5,14,37.5,14</points>
<intersection>35.5 0</intersection>
<intersection>37.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,13.5,16,15</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<connection>
<GID>65</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,13.5,17,15</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>15 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>17,15,18,15</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>19,13.5,22,13.5</points>
<connection>
<GID>66</GID>
<name>IN_3</name></connection>
<intersection>22 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22,13.5,22,15</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>13.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>20,14,20,15</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>18,14,20,14</points>
<intersection>18 3</intersection>
<intersection>20 1</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18,13.5,18,14</points>
<connection>
<GID>66</GID>
<name>IN_2</name></connection>
<intersection>14 2</intersection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>19,9,19,9.5</points>
<connection>
<GID>53</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>66</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>18,9,18,9.5</points>
<connection>
<GID>53</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>66</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>17,9,17,9.5</points>
<connection>
<GID>53</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>66</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>16,9,16,9.5</points>
<connection>
<GID>53</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,6,40.5,7</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,6,40.5,6</points>
<connection>
<GID>52</GID>
<name>carry_in</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,35,60.5,56</points>
<intersection>35 1</intersection>
<intersection>36 4</intersection>
<intersection>37 6</intersection>
<intersection>56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,35,71.5,35</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,56,60.5,56</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>60.5,36,71.5,36</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>60.5,37,61.5,37</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65.5,37,71.5,37</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,38,71.5,38</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,38,62,54</points>
<intersection>38 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,38,66,38</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,54,62,54</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61.5,39,71.5,39</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51,40,71.5,40</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-25,23.5,-25</points>
<connection>
<GID>96</GID>
<name>carry_in</name></connection>
<connection>
<GID>95</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-22,29.5,-21.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>31,-21.5,31,-21</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-21.5,31,-21.5</points>
<intersection>29.5 0</intersection>
<intersection>31 1</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-22,28.5,-21.5</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>29,-21.5,29,-21</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-21.5,29,-21.5</points>
<intersection>28.5 0</intersection>
<intersection>29 1</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-22,27.5,-21.5</points>
<connection>
<GID>95</GID>
<name>IN_2</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>27,-21.5,27,-21</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27,-21.5,27.5,-21.5</points>
<intersection>27 1</intersection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-21.5,25,-21</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>26.5,-22,26.5,-21.5</points>
<connection>
<GID>95</GID>
<name>IN_3</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>25,-21.5,26.5,-21.5</points>
<intersection>25 0</intersection>
<intersection>26.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-22,12,-21.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>13,-21.5,13,-21</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>12,-21.5,13,-21.5</points>
<intersection>12 0</intersection>
<intersection>13 1</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-22,11,-21</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<connection>
<GID>88</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-22,10,-21</points>
<connection>
<GID>96</GID>
<name>IN_2</name></connection>
<intersection>-21 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>9,-21,10,-21</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-22,7,-21</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>7,-22,9,-22</points>
<connection>
<GID>96</GID>
<name>IN_3</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>33,-41,33,-30</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-25,40.5,-25</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<connection>
<GID>95</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>4.5,-27,6,-27</points>
<connection>
<GID>96</GID>
<name>overflow</name></connection>
<intersection>4.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>4.5,-31,4.5,-27</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>-27 2</intersection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>36.5,-22,37.5,-22</points>
<connection>
<GID>95</GID>
<name>IN_B_0</name></connection>
<intersection>37.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>37.5,-22,37.5,-21</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<intersection>-22 0</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-22,18,-21</points>
<connection>
<GID>96</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-21.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>18,-21.5,19,-21.5</points>
<intersection>18 0</intersection>
<intersection>19 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>19,-22,19,-21.5</points>
<connection>
<GID>96</GID>
<name>IN_B_0</name></connection>
<intersection>-21.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-22,33.5,-21</points>
<connection>
<GID>95</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>-21.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>33.5,-21.5,35.5,-21.5</points>
<intersection>33.5 0</intersection>
<intersection>34.5 5</intersection>
<intersection>35.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>35.5,-22,35.5,-21.5</points>
<connection>
<GID>95</GID>
<name>IN_B_1</name></connection>
<intersection>-21.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>34.5,-22,34.5,-21.5</points>
<connection>
<GID>95</GID>
<name>IN_B_2</name></connection>
<intersection>-21.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-30,32,-30</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<connection>
<GID>95</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-41,31,-30</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<connection>
<GID>95</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-30,30,-30</points>
<connection>
<GID>95</GID>
<name>OUT_3</name></connection>
<connection>
<GID>105</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-30,15.5,-30</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<connection>
<GID>106</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-41,14.5,-30</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<connection>
<GID>96</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-30,13.5,-30</points>
<connection>
<GID>96</GID>
<name>OUT_2</name></connection>
<connection>
<GID>108</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-41,12.5,-30</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<connection>
<GID>96</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61.5,41.5,71.5,41.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>71.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71.5,41,71.5,42</points>
<connection>
<GID>8</GID>
<name>IN_7</name></connection>
<connection>
<GID>8</GID>
<name>IN_6</name></connection>
<intersection>41.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,42.5,-22.5,42.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<connection>
<GID>111</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,44.5,-22.5,44.5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<connection>
<GID>111</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,43.5,-16.5,43.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<connection>
<GID>111</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,38.5,-22.5,38.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<connection>
<GID>117</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,40.5,-22.5,40.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<connection>
<GID>117</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,39.5,-16.5,39.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<connection>
<GID>117</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,34.5,-22.5,34.5</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<connection>
<GID>125</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,36.5,-22.5,36.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<connection>
<GID>125</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,35.5,-16.5,35.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<connection>
<GID>125</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,30.5,-22.5,30.5</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<connection>
<GID>133</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,32.5,-22.5,32.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,31.5,-16.5,31.5</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<connection>
<GID>133</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,26.5,-22.5,26.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<connection>
<GID>141</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,28.5,-22.5,28.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<connection>
<GID>141</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,27.5,-16.5,27.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<connection>
<GID>141</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,22.5,-22.5,22.5</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<connection>
<GID>149</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,24.5,-22.5,24.5</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<connection>
<GID>149</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,23.5,-16.5,23.5</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<connection>
<GID>149</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,18.5,-22.5,18.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<connection>
<GID>157</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,20.5,-22.5,20.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<connection>
<GID>157</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,19.5,-16.5,19.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<connection>
<GID>157</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,14.5,-22.5,14.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<connection>
<GID>164</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,16.5,-22.5,16.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<connection>
<GID>164</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,15.5,-16.5,15.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<connection>
<GID>164</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,6.5,-22.5,6.5</points>
<connection>
<GID>193</GID>
<name>IN_1</name></connection>
<connection>
<GID>173</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,8.5,-22.5,8.5</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<connection>
<GID>172</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,4.5,-22.5,4.5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<connection>
<GID>175</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,2.5,-22.5,2.5</points>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<connection>
<GID>176</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-1.5,-22.5,-1.5</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<connection>
<GID>181</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,0.5,-22.5,0.5</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<connection>
<GID>179</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-3.5,-22.5,-3.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<connection>
<GID>182</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-5.5,-22.5,-5.5</points>
<connection>
<GID>196</GID>
<name>IN_1</name></connection>
<connection>
<GID>184</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-7.5,-22.5,-7.5</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<connection>
<GID>170</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-9.5,-22.5,-9.5</points>
<connection>
<GID>197</GID>
<name>IN_1</name></connection>
<connection>
<GID>186</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-13.5,-22.5,-13.5</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<connection>
<GID>188</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-11.5,-22.5,-11.5</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<connection>
<GID>148</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-15.5,-22.5,-15.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-17.5,-22.5,-17.5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<connection>
<GID>190</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-19.5,-22.5,-19.5</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<connection>
<GID>163</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-21.5,-22.5,-21.5</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<connection>
<GID>192</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,7.5,-16.5,7.5</points>
<connection>
<GID>193</GID>
<name>OUT</name></connection>
<connection>
<GID>202</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,3.5,-16.5,3.5</points>
<connection>
<GID>195</GID>
<name>OUT</name></connection>
<connection>
<GID>203</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-0.5,-16.5,-0.5</points>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<connection>
<GID>204</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-4.5,-16.5,-4.5</points>
<connection>
<GID>196</GID>
<name>OUT</name></connection>
<connection>
<GID>205</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-8.5,-16.5,-8.5</points>
<connection>
<GID>197</GID>
<name>OUT</name></connection>
<connection>
<GID>207</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-12.5,-16.5,-12.5</points>
<connection>
<GID>199</GID>
<name>OUT</name></connection>
<connection>
<GID>77</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-16.5,-16.5,-16.5</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<connection>
<GID>208</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-20.5,-16.5,-20.5</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<connection>
<GID>209</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-25.5,-22.5,-25.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<connection>
<GID>213</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-27.5,-22.5,-27.5</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<connection>
<GID>214</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-35.5,-22.5,-35.5</points>
<connection>
<GID>223</GID>
<name>IN_1</name></connection>
<connection>
<GID>84</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-33.5,-22.5,-33.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<connection>
<GID>216</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-37.5,-22.5,-37.5</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<connection>
<GID>217</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-39.5,-22.5,-39.5</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<connection>
<GID>80</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-43.5,-22.5,-43.5</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<connection>
<GID>218</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-41.5,-22.5,-41.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<connection>
<GID>212</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-47.5,-22.5,-47.5</points>
<connection>
<GID>226</GID>
<name>IN_1</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-45.5,-22.5,-45.5</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<connection>
<GID>210</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-51.5,-22.5,-51.5</points>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<connection>
<GID>219</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-49.5,-22.5,-49.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<connection>
<GID>90</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-55.5,-22.5,-55.5</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<connection>
<GID>228</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-53.5,-22.5,-53.5</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<connection>
<GID>228</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-29.5,-22.5,-29.5</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<connection>
<GID>82</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-31.5,-22.5,-31.5</points>
<connection>
<GID>222</GID>
<name>IN_1</name></connection>
<connection>
<GID>215</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-26.5,-16.5,-26.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<connection>
<GID>221</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-30.5,-16.5,-30.5</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<connection>
<GID>222</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-34.5,-16.5,-34.5</points>
<connection>
<GID>223</GID>
<name>OUT</name></connection>
<connection>
<GID>231</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-38.5,-16.5,-38.5</points>
<connection>
<GID>224</GID>
<name>OUT</name></connection>
<connection>
<GID>232</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-42.5,-16.5,-42.5</points>
<connection>
<GID>225</GID>
<name>OUT</name></connection>
<connection>
<GID>233</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-46.5,-16.5,-46.5</points>
<connection>
<GID>226</GID>
<name>OUT</name></connection>
<connection>
<GID>235</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-50.5,-16.5,-50.5</points>
<connection>
<GID>227</GID>
<name>OUT</name></connection>
<connection>
<GID>236</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-54.5,-16.5,-54.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<connection>
<GID>228</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>71,43,71.5,43</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,44,71.5,44</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>71,45,71.5,45</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-71.5,12.5,-71.5</points>
<connection>
<GID>242</GID>
<name>in_A_greater_B</name></connection>
<connection>
<GID>115</GID>
<name>A_greater_B</name></connection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-75.5,12.5,-75.5</points>
<connection>
<GID>242</GID>
<name>in_A_less_B</name></connection>
<connection>
<GID>115</GID>
<name>A_less_B</name></connection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-73.5,12.5,-73.5</points>
<connection>
<GID>242</GID>
<name>in_A_equal_B</name></connection>
<connection>
<GID>115</GID>
<name>A_equal_B</name></connection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-69.5,18.5,-69.5</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<connection>
<GID>115</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-69.5,16.5,-69.5</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<connection>
<GID>115</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-69.5,23.5,-69.5</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<connection>
<GID>115</GID>
<name>IN_B_2</name></connection></vsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-69.5,25.5,-69.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<connection>
<GID>115</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-69.5,24.5,-64.5</points>
<connection>
<GID>115</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>253</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-69.5,22.5,-64.5</points>
<connection>
<GID>115</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>243</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-69.5,17.5,-64.5</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<connection>
<GID>140</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-69.5,15.5,-64.5</points>
<connection>
<GID>115</GID>
<name>IN_3</name></connection>
<connection>
<GID>254</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-69.5,7,-69.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<connection>
<GID>242</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-69.5,5,-69.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<connection>
<GID>242</GID>
<name>IN_B_2</name></connection></vsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-69.5,6,-64.5</points>
<connection>
<GID>242</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>128</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-69.5,4,-64.5</points>
<connection>
<GID>242</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>152</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.38498e-008,-69.5,2.38498e-008,-69.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<connection>
<GID>242</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-69.5,-2,-69.5</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<connection>
<GID>242</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-69.5,-3,-64.5</points>
<connection>
<GID>242</GID>
<name>IN_3</name></connection>
<connection>
<GID>250</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-69.5,-1,-64.5</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<connection>
<GID>248</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-76.5,-6,-75.5</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<connection>
<GID>242</GID>
<name>A_less_B</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-76.5,-6,-76.5</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16,-73.5,-6,-73.5</points>
<connection>
<GID>242</GID>
<name>A_equal_B</name></connection>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>-16 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-16,-74.5,-16,-72.5</points>
<connection>
<GID>263</GID>
<name>IN_1</name></connection>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>-73.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-71.5,-6,-70.5</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<connection>
<GID>242</GID>
<name>A_greater_B</name></connection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-70.5,-6,-70.5</points>
<connection>
<GID>262</GID>
<name>IN_1</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-71.5,-22,-71.5</points>
<connection>
<GID>262</GID>
<name>OUT</name></connection>
<connection>
<GID>265</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-75.5,-22,-75.5</points>
<connection>
<GID>263</GID>
<name>OUT</name></connection>
<connection>
<GID>266</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,50,71.5,50</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>71,49,71.5,49</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>71,47,71.5,47</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,48,71.5,48</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,46,71.5,46</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>77.5,8,78,8</points>
<connection>
<GID>279</GID>
<name>OUT</name></connection>
<connection>
<GID>278</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>74,17.5,74,18.5</points>
<connection>
<GID>279</GID>
<name>SEL_2</name></connection>
<connection>
<GID>283</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,17.5,73,23.5</points>
<connection>
<GID>279</GID>
<name>SEL_3</name></connection>
<connection>
<GID>284</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,17.5,75,23.5</points>
<connection>
<GID>279</GID>
<name>SEL_1</name></connection>
<connection>
<GID>282</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>76,17.5,76,18.5</points>
<connection>
<GID>279</GID>
<name>SEL_0</name></connection>
<connection>
<GID>281</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,0.5,60.5,21.5</points>
<intersection>0.5 1</intersection>
<intersection>1.5 4</intersection>
<intersection>2.5 6</intersection>
<intersection>21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,0.5,71.5,0.5</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,21.5,60.5,21.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>60.5,1.5,71.5,1.5</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>60.5,2.5,61.5,2.5</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65.5,2.5,71.5,2.5</points>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,3.5,71.5,3.5</points>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,3.5,62,19.5</points>
<intersection>3.5 1</intersection>
<intersection>19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,3.5,66,3.5</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,19.5,62,19.5</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61.5,4.5,71.5,4.5</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51,5.5,71.5,5.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61.5,7,71.5,7</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>71.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71.5,6.5,71.5,7.5</points>
<connection>
<GID>279</GID>
<name>IN_7</name></connection>
<connection>
<GID>279</GID>
<name>IN_6</name></connection>
<intersection>7 1</intersection></vsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,8.5,71.5,8.5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,9.5,71.5,9.5</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,10.5,71.5,10.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,15.5,71.5,15.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,14.5,71.5,14.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,12.5,71.5,12.5</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,13.5,71.5,13.5</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,11.5,71.5,11.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>76.5,-29,77,-29</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<connection>
<GID>301</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-19.5,73,-18.5</points>
<connection>
<GID>302</GID>
<name>SEL_2</name></connection>
<connection>
<GID>4</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-19.5,72,-13.5</points>
<connection>
<GID>302</GID>
<name>SEL_3</name></connection>
<connection>
<GID>307</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-19.5,74,-13.5</points>
<connection>
<GID>302</GID>
<name>SEL_1</name></connection>
<connection>
<GID>305</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-19.5,75,-18.5</points>
<connection>
<GID>302</GID>
<name>SEL_0</name></connection>
<connection>
<GID>17</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-36.5,59.5,-15.5</points>
<intersection>-36.5 1</intersection>
<intersection>-35.5 4</intersection>
<intersection>-34.5 7</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-36.5,70.5,-36.5</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-15.5,59.5,-15.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>59.5,-35.5,70.5,-35.5</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>59.5,-34.5,60.5,-34.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-34.5,70.5,-34.5</points>
<connection>
<GID>308</GID>
<name>OUT_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69,-33.5,70.5,-33.5</points>
<connection>
<GID>309</GID>
<name>OUT_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-33.5,61,-17.5</points>
<intersection>-33.5 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-33.5,65,-33.5</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-17.5,61,-17.5</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-32.5,70.5,-32.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-31.5,70.5,-31.5</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-30,70.5,-30</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>70.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>70.5,-30.5,70.5,-29.5</points>
<connection>
<GID>302</GID>
<name>IN_7</name></connection>
<connection>
<GID>302</GID>
<name>IN_6</name></connection>
<intersection>-30 1</intersection></vsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-28.5,70.5,-28.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-27.5,70.5,-27.5</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>70,-26.5,70.5,-26.5</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-21.5,70.5,-21.5</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>70,-22.5,70.5,-22.5</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-24.5,70.5,-24.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-23.5,70.5,-23.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-25.5,70.5,-25.5</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76.5,-64.5,77,-64.5</points>
<connection>
<GID>318</GID>
<name>OUT</name></connection>
<connection>
<GID>238</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>73,-55,73,-54</points>
<connection>
<GID>318</GID>
<name>SEL_2</name></connection>
<connection>
<GID>320</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-55,72,-49</points>
<connection>
<GID>318</GID>
<name>SEL_3</name></connection>
<connection>
<GID>306</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-55,74,-49</points>
<connection>
<GID>318</GID>
<name>SEL_1</name></connection>
<connection>
<GID>118</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>75,-55,75,-54</points>
<connection>
<GID>318</GID>
<name>SEL_0</name></connection>
<connection>
<GID>319</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-72,59.5,-51</points>
<intersection>-72 1</intersection>
<intersection>-71 4</intersection>
<intersection>-70 7</intersection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-72,70.5,-72</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-51,59.5,-51</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>59.5,-71,70.5,-71</points>
<connection>
<GID>318</GID>
<name>IN_1</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>59.5,-70,60.5,-70</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-70,70.5,-70</points>
<connection>
<GID>321</GID>
<name>OUT_0</name></connection>
<connection>
<GID>318</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69,-69,70.5,-69</points>
<connection>
<GID>322</GID>
<name>OUT_0</name></connection>
<connection>
<GID>318</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-69,61,-53</points>
<intersection>-69 1</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-69,65,-69</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-53,61,-53</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-68,70.5,-68</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<connection>
<GID>318</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-67,70.5,-67</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<connection>
<GID>318</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-65.5,70.5,-65.5</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>70.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>70.5,-66,70.5,-65</points>
<connection>
<GID>318</GID>
<name>IN_7</name></connection>
<connection>
<GID>318</GID>
<name>IN_6</name></connection>
<intersection>-65.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-64,70.5,-64</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<connection>
<GID>318</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-63,70.5,-63</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<connection>
<GID>318</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-62,70.5,-62</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<connection>
<GID>318</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-57,70.5,-57</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<connection>
<GID>318</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-58,70.5,-58</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<connection>
<GID>318</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-60,70.5,-60</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<connection>
<GID>318</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-59,70.5,-59</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<connection>
<GID>318</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-61,70.5,-61</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<connection>
<GID>318</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121,42.5,121.5,42.5</points>
<connection>
<GID>331</GID>
<name>OUT</name></connection>
<connection>
<GID>329</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>117.5,52,117.5,53</points>
<connection>
<GID>331</GID>
<name>SEL_2</name></connection>
<connection>
<GID>333</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,52,116.5,58</points>
<connection>
<GID>331</GID>
<name>SEL_3</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,52,118.5,58</points>
<connection>
<GID>331</GID>
<name>SEL_1</name></connection>
<connection>
<GID>267</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,52,119.5,53</points>
<connection>
<GID>331</GID>
<name>SEL_0</name></connection>
<connection>
<GID>139</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,35,104,56</points>
<intersection>35 1</intersection>
<intersection>36 4</intersection>
<intersection>37 6</intersection>
<intersection>56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,35,115,35</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94,56,104,56</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>104,36,115,36</points>
<connection>
<GID>331</GID>
<name>IN_1</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>104,37,105,37</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,37,115,37</points>
<connection>
<GID>334</GID>
<name>OUT_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>113.5,38,115,38</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,38,105.5,54</points>
<intersection>38 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,38,109.5,38</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94,54,105.5,54</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,39,115,39</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94.5,40,115,40</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,41.5,115,41.5</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>115 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>115,41,115,42</points>
<connection>
<GID>331</GID>
<name>IN_7</name></connection>
<connection>
<GID>331</GID>
<name>IN_6</name></connection>
<intersection>41.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>114.5,43,115,43</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,44,115,44</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>114.5,45,115,45</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,50,115,50</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>114.5,49,115,49</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>114.5,47,115,47</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,48,115,48</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,46,115,46</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>121,8,121.5,8</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<connection>
<GID>341</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>117.5,17.5,117.5,18.5</points>
<connection>
<GID>162</GID>
<name>SEL_2</name></connection>
<connection>
<GID>269</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>116.5,17.5,116.5,23.5</points>
<connection>
<GID>162</GID>
<name>SEL_3</name></connection>
<connection>
<GID>343</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>118.5,17.5,118.5,23.5</points>
<connection>
<GID>162</GID>
<name>SEL_1</name></connection>
<connection>
<GID>244</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>119.5,17.5,119.5,18.5</points>
<connection>
<GID>162</GID>
<name>SEL_0</name></connection>
<connection>
<GID>342</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,0.5,104,21.5</points>
<intersection>0.5 1</intersection>
<intersection>1.5 4</intersection>
<intersection>2.5 6</intersection>
<intersection>21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,0.5,115,0.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94,21.5,104,21.5</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>104,1.5,115,1.5</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>104,2.5,105,2.5</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,2.5,115,2.5</points>
<connection>
<GID>249</GID>
<name>OUT_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,3.5,115,3.5</points>
<connection>
<GID>273</GID>
<name>OUT_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,3.5,105.5,19.5</points>
<intersection>3.5 1</intersection>
<intersection>19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,3.5,109.5,3.5</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94,19.5,105.5,19.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,4.5,115,4.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94.5,5.5,115,5.5</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,7,115,7</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>115 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>115,6.5,115,7.5</points>
<connection>
<GID>162</GID>
<name>IN_7</name></connection>
<connection>
<GID>162</GID>
<name>IN_6</name></connection>
<intersection>7 1</intersection></vsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114.5,8.5,115,8.5</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,9.5,115,9.5</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114.5,10.5,115,10.5</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,15.5,115,15.5</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114.5,14.5,115,14.5</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114.5,12.5,115,12.5</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,13.5,115,13.5</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,11.5,115,11.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>120,-29,120.5,-29</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<connection>
<GID>355</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>116.5,-19.5,116.5,-18.5</points>
<connection>
<GID>187</GID>
<name>SEL_2</name></connection>
<connection>
<GID>261</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>115.5,-19.5,115.5,-13.5</points>
<connection>
<GID>187</GID>
<name>SEL_3</name></connection>
<connection>
<GID>359</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>117.5,-19.5,117.5,-13.5</points>
<connection>
<GID>187</GID>
<name>SEL_1</name></connection>
<connection>
<GID>358</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>118.5,-19.5,118.5,-18.5</points>
<connection>
<GID>187</GID>
<name>SEL_0</name></connection>
<connection>
<GID>247</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-36.5,103,-15.5</points>
<intersection>-36.5 1</intersection>
<intersection>-35.5 4</intersection>
<intersection>-34.5 7</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103,-36.5,114,-36.5</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93,-15.5,103,-15.5</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>103,-35.5,114,-35.5</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>103,-34.5,104,-34.5</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-34.5,114,-34.5</points>
<connection>
<GID>360</GID>
<name>OUT_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>112.5,-33.5,114,-33.5</points>
<connection>
<GID>361</GID>
<name>OUT_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-33.5,104.5,-17.5</points>
<intersection>-33.5 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-33.5,108.5,-33.5</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93,-17.5,104.5,-17.5</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-32.5,114,-32.5</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,-31.5,114,-31.5</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-30,114,-30</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>114 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114,-30.5,114,-29.5</points>
<connection>
<GID>187</GID>
<name>IN_7</name></connection>
<connection>
<GID>187</GID>
<name>IN_6</name></connection>
<intersection>-30 1</intersection></vsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>113.5,-28.5,114,-28.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-27.5,114,-27.5</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>113.5,-26.5,114,-26.5</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-21.5,114,-21.5</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>113.5,-22.5,114,-22.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-24.5,114,-24.5</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-23.5,114,-23.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-25.5,114,-25.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-64.5,120.5,-64.5</points>
<connection>
<GID>367</GID>
<name>OUT</name></connection>
<connection>
<GID>158</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>116.5,-55,116.5,-54</points>
<connection>
<GID>367</GID>
<name>SEL_2</name></connection>
<connection>
<GID>368</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-55,115.5,-49</points>
<connection>
<GID>367</GID>
<name>SEL_3</name></connection>
<connection>
<GID>189</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-55,117.5,-49</points>
<connection>
<GID>367</GID>
<name>SEL_1</name></connection>
<connection>
<GID>150</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-55,118.5,-54</points>
<connection>
<GID>367</GID>
<name>SEL_0</name></connection>
<connection>
<GID>198</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-72,103,-51</points>
<intersection>-72 1</intersection>
<intersection>-71 4</intersection>
<intersection>-70 7</intersection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103,-72,114,-72</points>
<connection>
<GID>367</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93,-51,103,-51</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>103,-71,114,-71</points>
<connection>
<GID>367</GID>
<name>IN_1</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>103,-70,104,-70</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-70,114,-70</points>
<connection>
<GID>369</GID>
<name>OUT_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>112.5,-69,114,-69</points>
<connection>
<GID>370</GID>
<name>OUT_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-69,104.5,-53</points>
<intersection>-69 1</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-69,108.5,-69</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93,-53,104.5,-53</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-68,114,-68</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,-67,114,-67</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-65.5,114,-65.5</points>
<connection>
<GID>371</GID>
<name>IN_0</name></connection>
<intersection>114 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114,-66,114,-65</points>
<connection>
<GID>367</GID>
<name>IN_7</name></connection>
<connection>
<GID>367</GID>
<name>IN_6</name></connection>
<intersection>-65.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>113.5,-64,114,-64</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-63,114,-63</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>113.5,-62,114,-62</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-57,114,-57</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>113.5,-58,114,-58</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-60,114,-60</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-59,114,-59</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-61,114,-61</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_11</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,44.2,-46.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,44.2,-46.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,44.2,-46.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,44.2,-46.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,44.2,-46.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,44.2,-46.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,44.2,-46.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,44.2,-46.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,44.2,-46.2</PageViewport></page 9></circuit>