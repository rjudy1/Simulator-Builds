
<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-32.95,39.6893,61.95,-63.2229</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>14.5,-13</position>
<gparam>LABEL_TEXT Go to https://cedar.to/vjyQw7 to download the latest version!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>14.5,-9.5</position>
<gparam>LABEL_TEXT Error: This file was made with a newer version of Cedar Logic!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate></page 0>
</circuit>
<throw_away></throw_away>

	<version>2.3.5 | 2018-09-25 23:06:05</version><circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0.968155,131.511,442.671,-84.5946</PageViewport>
<gate>
<ID>65</ID>
<type>DA_FROM</type>
<position>27.5,78.5</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID vdd</lparam></gate>
<gate>
<ID>1</ID>
<type>DA_FROM</type>
<position>28.5,71.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir12</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_AND2</type>
<position>125.5,-42</position>
<input>
<ID>IN_0</ID>316 </input>
<input>
<ID>IN_1</ID>317 </input>
<output>
<ID>OUT</ID>321 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>104,159</position>
<gparam>LABEL_TEXT MANO MACHINE CCL</gparam>
<gparam>TEXT_HEIGHT 8</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>3</ID>
<type>DA_FROM</type>
<position>49.5,-19</position>
<input>
<ID>IN_0</ID>296 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr12</lparam></gate>
<gate>
<ID>4</ID>
<type>DA_FROM</type>
<position>18,74</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir14</lparam></gate>
<gate>
<ID>5</ID>
<type>DE_TO</type>
<position>145,25</position>
<input>
<ID>IN_0</ID>315 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcBus</lparam></gate>
<gate>
<ID>6</ID>
<type>EE_VDD</type>
<position>-42,18.5</position>
<output>
<ID>OUT_0</ID>351 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>7</ID>
<type>DA_FROM</type>
<position>118,-23.5</position>
<input>
<ID>IN_0</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>8</ID>
<type>DA_FROM</type>
<position>54.5,130.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID vdd</lparam></gate>
<gate>
<ID>10</ID>
<type>DE_TO</type>
<position>46,82</position>
<input>
<ID>IN_0</ID>38 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D7</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>134.5,32.5</position>
<gparam>LABEL_TEXT PC Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>DE_TO</type>
<position>77.5,118.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_AND3</type>
<position>-72,11</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>269 </input>
<input>
<ID>IN_2</ID>270 </input>
<output>
<ID>OUT</ID>339 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>16</ID>
<type>DE_TO</type>
<position>77,122.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T7</lparam></gate>
<gate>
<ID>17</ID>
<type>DA_FROM</type>
<position>53.5,-7</position>
<input>
<ID>IN_0</ID>285 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr1</lparam></gate>
<gate>
<ID>19</ID>
<type>DA_FROM</type>
<position>-81,-11.5</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir7</lparam></gate>
<gate>
<ID>20</ID>
<type>DE_TO</type>
<position>81.5,115.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>-17,112</position>
<input>
<ID>IN_0</ID>196 </input>
<input>
<ID>IN_1</ID>195 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>DA_FROM</type>
<position>45.5,121.5</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>391</ID>
<type>DA_FROM</type>
<position>-81,11</position>
<input>
<ID>IN_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir6</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>47,-12</position>
<input>
<ID>IN_0</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr6</lparam></gate>
<gate>
<ID>25</ID>
<type>DE_TO</type>
<position>77,130.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T15</lparam></gate>
<gate>
<ID>385</ID>
<type>AE_OR3</type>
<position>144.5,100.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>56 </input>
<input>
<ID>IN_2</ID>61 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_AND2</type>
<position>39,56</position>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>204 </input>
<output>
<ID>OUT</ID>255 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>DE_TO</type>
<position>81.5,127.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T12</lparam></gate>
<gate>
<ID>28</ID>
<type>DA_FROM</type>
<position>118.5,-48.5</position>
<input>
<ID>IN_0</ID>319 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>389</ID>
<type>DE_TO</type>
<position>53.5,56</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /I</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>-81,-18</position>
<input>
<ID>IN_0</ID>333 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir6</lparam></gate>
<gate>
<ID>399</ID>
<type>DA_FROM</type>
<position>195.5,-12</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>51,-17.5</position>
<input>
<ID>IN_0</ID>295 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr11</lparam></gate>
<gate>
<ID>33</ID>
<type>DE_TO</type>
<position>77,124.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T9</lparam></gate>
<gate>
<ID>393</ID>
<type>DA_FROM</type>
<position>122.5,136</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>-22,111</position>
<input>
<ID>IN_0</ID>195 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>44,124</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>-15,95</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>387</ID>
<type>AA_AND2</type>
<position>131.5,137</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>DE_TO</type>
<position>78,116.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>397</ID>
<type>DA_FROM</type>
<position>115,119</position>
<input>
<ID>IN_0</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>38</ID>
<type>DA_FROM</type>
<position>-81,9</position>
<input>
<ID>IN_0</ID>270 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>39</ID>
<type>BI_DECODER_4x16</type>
<position>61.5,123</position>
<input>
<ID>ENABLE</ID>12 </input>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>22 </input>
<input>
<ID>IN_2</ID>21 </input>
<input>
<ID>IN_3</ID>23 </input>
<output>
<ID>OUT_0</ID>18 </output>
<output>
<ID>OUT_1</ID>17 </output>
<output>
<ID>OUT_10</ID>6 </output>
<output>
<ID>OUT_11</ID>5 </output>
<output>
<ID>OUT_12</ID>4 </output>
<output>
<ID>OUT_13</ID>3 </output>
<output>
<ID>OUT_14</ID>2 </output>
<output>
<ID>OUT_15</ID>1 </output>
<output>
<ID>OUT_2</ID>16 </output>
<output>
<ID>OUT_3</ID>15 </output>
<output>
<ID>OUT_4</ID>14 </output>
<output>
<ID>OUT_5</ID>13 </output>
<output>
<ID>OUT_6</ID>10 </output>
<output>
<ID>OUT_7</ID>9 </output>
<output>
<ID>OUT_8</ID>8 </output>
<output>
<ID>OUT_9</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>407</ID>
<type>DA_FROM</type>
<position>75,61</position>
<input>
<ID>IN_0</ID>205 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID start</lparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>80.5,-15</position>
<input>
<ID>IN_0</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID zeroDR</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_REGISTER4</type>
<position>48.5,116.5</position>
<output>
<ID>OUT_0</ID>24 </output>
<output>
<ID>OUT_1</ID>22 </output>
<output>
<ID>OUT_2</ID>21 </output>
<output>
<ID>OUT_3</ID>23 </output>
<input>
<ID>clear</ID>28 </input>
<input>
<ID>clock</ID>25 </input>
<input>
<ID>count_enable</ID>26 </input>
<input>
<ID>load</ID>27 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>401</ID>
<type>FF_GND</type>
<position>209.5,-26.5</position>
<output>
<ID>OUT_0</ID>174 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>AE_OR4</type>
<position>8,115.5</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>202 </input>
<input>
<ID>IN_2</ID>203 </input>
<input>
<ID>IN_3</ID>1194 </input>
<output>
<ID>OUT</ID>180 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>43</ID>
<type>DA_FROM</type>
<position>42.5,112</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>395</ID>
<type>DA_FROM</type>
<position>115,123</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>44</ID>
<type>DA_FROM</type>
<position>-82,45.5</position>
<input>
<ID>IN_0</ID>323 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID start</lparam></gate>
<gate>
<ID>45</ID>
<type>DA_FROM</type>
<position>42.5,109</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrSC</lparam></gate>
<gate>
<ID>405</ID>
<type>DA_FROM</type>
<position>79,63</position>
<input>
<ID>IN_0</ID>188 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_AND2</type>
<position>29.5,61.5</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>251 </input>
<output>
<ID>OUT</ID>252 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>81.5,129.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T14</lparam></gate>
<gate>
<ID>415</ID>
<type>DA_FROM</type>
<position>120,-32.5</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_AND3</type>
<position>125.5,-13</position>
<input>
<ID>IN_0</ID>303 </input>
<input>
<ID>IN_1</ID>302 </input>
<input>
<ID>IN_2</ID>304 </input>
<output>
<ID>OUT</ID>305 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>49</ID>
<type>DE_TO</type>
<position>77,128.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T13</lparam></gate>
<gate>
<ID>409</ID>
<type>DE_TO</type>
<position>92,57</position>
<input>
<ID>IN_0</ID>232 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incTR</lparam></gate>
<gate>
<ID>50</ID>
<type>DE_TO</type>
<position>77,126.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T11</lparam></gate>
<gate>
<ID>51</ID>
<type>DA_FROM</type>
<position>120,-28.5</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGO</lparam></gate>
<gate>
<ID>403</ID>
<type>AA_AND2</type>
<position>85,64</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>DE_TO</type>
<position>82,125.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T10</lparam></gate>
<gate>
<ID>53</ID>
<type>DA_FROM</type>
<position>120,18.5</position>
<input>
<ID>IN_0</ID>274 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>413</ID>
<type>AA_AND2</type>
<position>125,-31.5</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>DE_TO</type>
<position>82,123.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T8</lparam></gate>
<gate>
<ID>55</ID>
<type>DE_TO</type>
<position>82,121.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>56</ID>
<type>DA_FROM</type>
<position>-5.5,22</position>
<input>
<ID>IN_0</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>423</ID>
<type>AA_AND2</type>
<position>-72,-23.5</position>
<input>
<ID>IN_0</ID>334 </input>
<input>
<ID>IN_1</ID>335 </input>
<output>
<ID>OUT</ID>344 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>DE_TO</type>
<position>77,120.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>58</ID>
<type>DE_TO</type>
<position>143,-55.5</position>
<input>
<ID>IN_0</ID>329 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrPC</lparam></gate>
<gate>
<ID>417</ID>
<type>DA_FROM</type>
<position>-48,12</position>
<input>
<ID>IN_0</ID>347 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>59</ID>
<type>DE_TO</type>
<position>82,119.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>60</ID>
<type>DE_TO</type>
<position>81.5,117.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>411</ID>
<type>AA_AND2</type>
<position>85,51.5</position>
<input>
<ID>IN_0</ID>234 </input>
<input>
<ID>IN_1</ID>250 </input>
<output>
<ID>OUT</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>AE_SMALL_INVERTER</type>
<position>41,82</position>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_OR4</type>
<position>-56,23.5</position>
<input>
<ID>IN_0</ID>336 </input>
<input>
<ID>IN_1</ID>337 </input>
<input>
<ID>IN_2</ID>338 </input>
<input>
<ID>IN_3</ID>339 </input>
<output>
<ID>OUT</ID>345 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>421</ID>
<type>DA_FROM</type>
<position>-81,4.5</position>
<input>
<ID>IN_0</ID>271 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>63</ID>
<type>BE_DECODER_3x8</type>
<position>34.5,75</position>
<input>
<ID>ENABLE</ID>29 </input>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>31 </input>
<input>
<ID>IN_2</ID>32 </input>
<output>
<ID>OUT_0</ID>33 </output>
<output>
<ID>OUT_1</ID>41 </output>
<output>
<ID>OUT_2</ID>40 </output>
<output>
<ID>OUT_3</ID>39 </output>
<output>
<ID>OUT_4</ID>37 </output>
<output>
<ID>OUT_5</ID>36 </output>
<output>
<ID>OUT_6</ID>35 </output>
<output>
<ID>OUT_7</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>118,-43</position>
<input>
<ID>IN_0</ID>317 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>66</ID>
<type>DA_FROM</type>
<position>120.5,12.5</position>
<input>
<ID>IN_0</ID>277 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>67</ID>
<type>DE_TO</type>
<position>47,78.5</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>68</ID>
<type>DE_TO</type>
<position>52.5,77.5</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>69</ID>
<type>DA_FROM</type>
<position>120,16.5</position>
<input>
<ID>IN_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>70</ID>
<type>DE_TO</type>
<position>47,76.5</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>210,29</position>
<input>
<ID>IN_0</ID>377 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>72</ID>
<type>DE_TO</type>
<position>52.5,75.5</position>
<input>
<ID>IN_0</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>73</ID>
<type>DA_FROM</type>
<position>-5.5,12.5</position>
<input>
<ID>IN_0</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>74</ID>
<type>DE_TO</type>
<position>47,74.5</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>4.5,85</position>
<gparam>LABEL_TEXT Instruction Decoder</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>DA_FROM</type>
<position>-7.5,-8.5</position>
<input>
<ID>IN_0</ID>215 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir7</lparam></gate>
<gate>
<ID>77</ID>
<type>DE_TO</type>
<position>52.5,73.5</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>-82,54</position>
<input>
<ID>IN_0</ID>325 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>79</ID>
<type>DE_TO</type>
<position>47,72.5</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>45.5,-13.5</position>
<input>
<ID>IN_0</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr7</lparam></gate>
<gate>
<ID>81</ID>
<type>DE_TO</type>
<position>52.5,71.5</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>23,72.5</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir13</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>130.5,26.5</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>135.5,87.5</position>
<gparam>LABEL_TEXT AR Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>DE_TO</type>
<position>156,10</position>
<input>
<ID>IN_0</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incPC</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>206.5,1.5</position>
<gparam>LABEL_TEXT IR Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>DA_FROM</type>
<position>195.5,-6.5</position>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>88</ID>
<type>DE_TO</type>
<position>214,-5.5</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldIR</lparam></gate>
<gate>
<ID>455</ID>
<type>DE_TO</type>
<position>149,42</position>
<input>
<ID>IN_0</ID>382 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrAR</lparam></gate>
<gate>
<ID>89</ID>
<type>DE_TO</type>
<position>156,130.5</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID read_memory</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>133.5,142.5</position>
<gparam>LABEL_TEXT Memory Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>449</ID>
<type>AE_SMALL_INVERTER</type>
<position>-88,26.5</position>
<input>
<ID>IN_0</ID>261 </input>
<output>
<ID>OUT_0</ID>352 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>91</ID>
<type>DA_FROM</type>
<position>205,74.5</position>
<input>
<ID>IN_0</ID>44 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>92</ID>
<type>DA_FROM</type>
<position>205,76.5</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir11</lparam></gate>
<gate>
<ID>93</ID>
<type>AA_AND2</type>
<position>210,75.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>371 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>DE_TO</type>
<position>222,73.5</position>
<input>
<ID>IN_0</ID>1199 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrAC</lparam></gate>
<gate>
<ID>453</ID>
<type>AA_AND2</type>
<position>215,28</position>
<input>
<ID>IN_0</ID>377 </input>
<input>
<ID>IN_1</ID>376 </input>
<output>
<ID>OUT</ID>378 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>201.5,82</position>
<gparam>LABEL_TEXT AC Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>DE_TO</type>
<position>225.5,52</position>
<input>
<ID>IN_0</ID>1198 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldAC</lparam></gate>
<gate>
<ID>463</ID>
<type>AE_SMALL_INVERTER</type>
<position>129.5,73</position>
<input>
<ID>IN_0</ID>396 </input>
<output>
<ID>OUT_0</ID>395 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>97</ID>
<type>DE_TO</type>
<position>-60,101</position>
<input>
<ID>IN_0</ID>229 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /IEN</lparam></gate>
<gate>
<ID>98</ID>
<type>DA_FROM</type>
<position>198,67.5</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>457</ID>
<type>DA_FROM</type>
<position>127,71</position>
<input>
<ID>IN_0</ID>389 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID I</lparam></gate>
<gate>
<ID>99</ID>
<type>EE_VDD</type>
<position>-67,140.5</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>100</ID>
<type>DA_FROM</type>
<position>120.5,-13</position>
<input>
<ID>IN_0</ID>302 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>451</ID>
<type>DA_FROM</type>
<position>211.5,72.5</position>
<input>
<ID>IN_0</ID>370 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID start</lparam></gate>
<gate>
<ID>101</ID>
<type>DE_TO</type>
<position>2,62</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>102</ID>
<type>DA_FROM</type>
<position>194.5,115.5</position>
<input>
<ID>IN_0</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>461</ID>
<type>DA_FROM</type>
<position>127.5,79.5</position>
<input>
<ID>IN_0</ID>386 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>103</ID>
<type>DE_TO</type>
<position>151,76</position>
<input>
<ID>IN_0</ID>391 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldAR</lparam></gate>
<gate>
<ID>104</ID>
<type>DA_FROM</type>
<position>198.5,65</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>105</ID>
<type>DA_FROM</type>
<position>198.5,63</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>106</ID>
<type>DA_FROM</type>
<position>127,75</position>
<input>
<ID>IN_0</ID>388 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>107</ID>
<type>DA_FROM</type>
<position>198.5,61</position>
<input>
<ID>IN_0</ID>53 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>108</ID>
<type>AE_OR3</type>
<position>203.5,63</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>53 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>459</ID>
<type>AA_AND2</type>
<position>135.5,80.5</position>
<input>
<ID>IN_0</ID>385 </input>
<input>
<ID>IN_1</ID>386 </input>
<output>
<ID>OUT</ID>392 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_AND2</type>
<position>211,65.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>168 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>DE_TO</type>
<position>220,28</position>
<input>
<ID>IN_0</ID>378 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incAC</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_AND3</type>
<position>135.5,71</position>
<input>
<ID>IN_0</ID>395 </input>
<input>
<ID>IN_1</ID>389 </input>
<input>
<ID>IN_2</ID>390 </input>
<output>
<ID>OUT</ID>394 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>112</ID>
<type>DA_FROM</type>
<position>206,51</position>
<input>
<ID>IN_0</ID>164 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>113</ID>
<type>DA_FROM</type>
<position>127,77</position>
<input>
<ID>IN_0</ID>387 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>114</ID>
<type>DA_FROM</type>
<position>198.5,47</position>
<input>
<ID>IN_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir6</lparam></gate>
<gate>
<ID>115</ID>
<type>DA_FROM</type>
<position>120.5,4.5</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir3</lparam></gate>
<gate>
<ID>116</ID>
<type>DA_FROM</type>
<position>120.5,10</position>
<input>
<ID>IN_0</ID>126 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir4</lparam></gate>
<gate>
<ID>117</ID>
<type>DA_FROM</type>
<position>120.5,-6</position>
<input>
<ID>IN_0</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /E</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_OR4</type>
<position>124.5,122</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>140 </input>
<input>
<ID>IN_2</ID>141 </input>
<input>
<ID>IN_3</ID>143 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_OR4</type>
<position>150,10</position>
<input>
<ID>IN_0</ID>276 </input>
<input>
<ID>IN_1</ID>279 </input>
<input>
<ID>IN_2</ID>305 </input>
<input>
<ID>IN_3</ID>105 </input>
<output>
<ID>OUT</ID>312 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>120</ID>
<type>DA_FROM</type>
<position>204.5,20.5</position>
<input>
<ID>IN_0</ID>171 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>121</ID>
<type>DA_FROM</type>
<position>-100.5,85</position>
<input>
<ID>IN_0</ID>231 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGO</lparam></gate>
<gate>
<ID>122</ID>
<type>DE_TO</type>
<position>223.5,15.5</position>
<input>
<ID>IN_0</ID>369 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acBus</lparam></gate>
<gate>
<ID>124</ID>
<type>DA_FROM</type>
<position>204.5,18.5</position>
<input>
<ID>IN_0</ID>172 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>195.5,-14</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>206,38</position>
<input>
<ID>IN_0</ID>166 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir11</lparam></gate>
<gate>
<ID>127</ID>
<type>DA_FROM</type>
<position>-81,32.5</position>
<input>
<ID>IN_0</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>-79,62</position>
<gparam>LABEL_TEXT Output Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>DA_FROM</type>
<position>206,55</position>
<input>
<ID>IN_0</ID>162 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>282</ID>
<type>AA_LABEL</type>
<position>-8,31.5</position>
<gparam>LABEL_TEXT ALU Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>DE_TO</type>
<position>-72,53</position>
<input>
<ID>IN_0</ID>324 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldOut</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>198.5,43</position>
<input>
<ID>IN_0</ID>159 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir9</lparam></gate>
<gate>
<ID>292</ID>
<type>AA_TOGGLE</type>
<position>-87.5,122</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>120.5,130.5</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID I</lparam></gate>
<gate>
<ID>133</ID>
<type>AE_OR2</type>
<position>216.5,73.5</position>
<input>
<ID>IN_0</ID>371 </input>
<input>
<ID>IN_1</ID>370 </input>
<output>
<ID>OUT</ID>1199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>286</ID>
<type>AA_TOGGLE</type>
<position>-86.5,137</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>134</ID>
<type>DA_FROM</type>
<position>-82,52</position>
<input>
<ID>IN_0</ID>326 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir10</lparam></gate>
<gate>
<ID>135</ID>
<type>DE_TO</type>
<position>151.5,100.5</position>
<input>
<ID>IN_0</ID>63 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID write_memory</lparam></gate>
<gate>
<ID>280</ID>
<type>AA_AND2</type>
<position>0,-14</position>
<input>
<ID>IN_0</ID>211 </input>
<input>
<ID>IN_1</ID>217 </input>
<output>
<ID>OUT</ID>218 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>DE_TO</type>
<position>14,115.5</position>
<input>
<ID>IN_0</ID>180 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrSC</lparam></gate>
<gate>
<ID>137</ID>
<type>DE_TO</type>
<position>143.5,63.5</position>
<input>
<ID>IN_0</ID>379 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incAR</lparam></gate>
<gate>
<ID>290</ID>
<type>DA_FROM</type>
<position>-89.5,134</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>138</ID>
<type>DE_TO</type>
<position>146.5,53.5</position>
<input>
<ID>IN_0</ID>357 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID arBus</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>203,133.5</position>
<gparam>LABEL_TEXT DR Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>300</ID>
<type>DE_TO</type>
<position>-59,137</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGI</lparam></gate>
<gate>
<ID>140</ID>
<type>DA_FROM</type>
<position>120,-18.5</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGI</lparam></gate>
<gate>
<ID>141</ID>
<type>DE_TO</type>
<position>215.5,121.5</position>
<input>
<ID>IN_0</ID>364 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldDR</lparam></gate>
<gate>
<ID>294</ID>
<type>BE_JKFF_LOW</type>
<position>-67,135</position>
<input>
<ID>J</ID>42 </input>
<input>
<ID>K</ID>67 </input>
<output>
<ID>Q</ID>62 </output>
<input>
<ID>clear</ID>1202 </input>
<input>
<ID>clock</ID>49 </input>
<output>
<ID>nQ</ID>66 </output>
<input>
<ID>set</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>988</ID>
<type>DA_FROM</type>
<position>-77.5,-27.5</position>
<input>
<ID>IN_0</ID>987 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID start</lparam></gate>
<gate>
<ID>142</ID>
<type>AE_OR3</type>
<position>133.5,-26.5</position>
<input>
<ID>IN_0</ID>1142 </input>
<input>
<ID>IN_1</ID>308 </input>
<input>
<ID>IN_2</ID>103 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>288</ID>
<type>DA_FROM</type>
<position>-90.5,119</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_AND2</type>
<position>208.5,121.5</position>
<input>
<ID>IN_0</ID>363 </input>
<input>
<ID>IN_1</ID>362 </input>
<output>
<ID>OUT</ID>364 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_AND2</type>
<position>137,107</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>298</ID>
<type>BE_JKFF_LOW</type>
<position>-67,120</position>
<input>
<ID>J</ID>46 </input>
<input>
<ID>K</ID>91 </input>
<output>
<ID>Q</ID>59 </output>
<input>
<ID>clear</ID>1202 </input>
<input>
<ID>clock</ID>57 </input>
<output>
<ID>nQ</ID>58 </output>
<input>
<ID>set</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>146</ID>
<type>DA_FROM</type>
<position>47,7.5</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>147</ID>
<type>AE_OR2</type>
<position>143.5,42</position>
<input>
<ID>IN_0</ID>383 </input>
<input>
<ID>IN_1</ID>384 </input>
<output>
<ID>OUT</ID>382 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>308</ID>
<type>DA_FROM</type>
<position>-15.5,64</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>148</ID>
<type>DE_OR8</type>
<position>62,1</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>77 </input>
<input>
<ID>IN_2</ID>78 </input>
<input>
<ID>IN_3</ID>79 </input>
<input>
<ID>IN_4</ID>83 </input>
<input>
<ID>IN_5</ID>82 </input>
<input>
<ID>IN_6</ID>81 </input>
<input>
<ID>IN_7</ID>80 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>996</ID>
<type>DA_FROM</type>
<position>120,-20.5</position>
<input>
<ID>IN_0</ID>306 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir9</lparam></gate>
<gate>
<ID>149</ID>
<type>DA_FROM</type>
<position>125.5,42</position>
<input>
<ID>IN_0</ID>381 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>302</ID>
<type>AA_AND2</type>
<position>-83,133</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>DA_FROM</type>
<position>48,-0.5</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>151</ID>
<type>DA_FROM</type>
<position>52,11.5</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>296</ID>
<type>DA_FROM</type>
<position>-74.5,135</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>152</ID>
<type>DE_OR8</type>
<position>62,10</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>69 </input>
<input>
<ID>IN_2</ID>70 </input>
<input>
<ID>IN_3</ID>71 </input>
<input>
<ID>IN_4</ID>75 </input>
<input>
<ID>IN_5</ID>74 </input>
<input>
<ID>IN_6</ID>73 </input>
<input>
<ID>IN_7</ID>72 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>153</ID>
<type>DA_FROM</type>
<position>127.5,81.5</position>
<input>
<ID>IN_0</ID>385 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>306</ID>
<type>AA_AND2</type>
<position>135.5,76</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>388 </input>
<output>
<ID>OUT</ID>393 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>154</ID>
<type>BE_NOR2</type>
<position>75,4.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>155</ID>
<type>DA_FROM</type>
<position>55.5,13.5</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>316</ID>
<type>AA_AND2</type>
<position>-78,81.5</position>
<input>
<ID>IN_0</ID>247 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>248 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>DA_FROM</type>
<position>53.5,12.5</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>157</ID>
<type>DA_FROM</type>
<position>51,10.5</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>310</ID>
<type>DA_FROM</type>
<position>-15.5,60</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>158</ID>
<type>DA_FROM</type>
<position>49.5,9.5</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>159</ID>
<type>DA_FROM</type>
<position>48,8.5</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>304</ID>
<type>AA_AND2</type>
<position>-84,118</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>160</ID>
<type>DA_FROM</type>
<position>45.5,6</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_AND2</type>
<position>-93.5,98</position>
<input>
<ID>IN_0</ID>224 </input>
<input>
<ID>IN_1</ID>225 </input>
<output>
<ID>OUT</ID>227 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>314</ID>
<type>DA_FROM</type>
<position>-15,54</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /I</lparam></gate>
<gate>
<ID>162</ID>
<type>DA_FROM</type>
<position>55.5,4.5</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>163</ID>
<type>DA_FROM</type>
<position>194.5,108</position>
<input>
<ID>IN_0</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>164</ID>
<type>DA_FROM</type>
<position>53.5,3.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_FROM</type>
<position>52,2.5</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>318</ID>
<type>BE_JKFF_LOW</type>
<position>70.5,97.5</position>
<input>
<ID>J</ID>175 </input>
<input>
<ID>K</ID>176 </input>
<output>
<ID>Q</ID>177 </output>
<input>
<ID>clear</ID>181 </input>
<input>
<ID>clock</ID>173 </input>
<output>
<ID>nQ</ID>178 </output>
<input>
<ID>set</ID>181 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>166</ID>
<type>AE_OR2</type>
<position>-95.5,86</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>231 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>167</ID>
<type>DA_FROM</type>
<position>51,1.5</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>312</ID>
<type>DE_TO</type>
<position>2.5,54</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>168</ID>
<type>DA_FROM</type>
<position>49.5,0.5</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>169</ID>
<type>DA_FROM</type>
<position>47,-1.5</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>170</ID>
<type>DA_FROM</type>
<position>46.5,-2.5</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>171</ID>
<type>DE_TO</type>
<position>81,4.5</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID zeroAC</lparam></gate>
<gate>
<ID>172</ID>
<type>DA_FROM</type>
<position>52,-16.5</position>
<input>
<ID>IN_0</ID>294 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr10</lparam></gate>
<gate>
<ID>173</ID>
<type>DA_FROM</type>
<position>48,-20</position>
<input>
<ID>IN_0</ID>297 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr13</lparam></gate>
<gate>
<ID>174</ID>
<type>DA_FROM</type>
<position>193.5,90.5</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID start</lparam></gate>
<gate>
<ID>175</ID>
<type>DA_FROM</type>
<position>128.5,109</position>
<input>
<ID>IN_0</ID>110 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>176</ID>
<type>DA_FROM</type>
<position>52,-8</position>
<input>
<ID>IN_0</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr2</lparam></gate>
<gate>
<ID>177</ID>
<type>DA_FROM</type>
<position>123,106</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>178</ID>
<type>DA_FROM</type>
<position>123,104</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>179</ID>
<type>AE_OR2</type>
<position>128,105</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>109 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>180</ID>
<type>AE_OR3</type>
<position>-11,103.5</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>145 </input>
<input>
<ID>IN_2</ID>151 </input>
<output>
<ID>OUT</ID>1193 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>181</ID>
<type>DA_FROM</type>
<position>48,-11</position>
<input>
<ID>IN_0</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr5</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_AND2</type>
<position>137,100.5</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_1</ID>113 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>183</ID>
<type>DE_TO</type>
<position>-59,84</position>
<input>
<ID>IN_0</ID>245 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>184</ID>
<type>DA_FROM</type>
<position>132,101.5</position>
<input>
<ID>IN_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>185</ID>
<type>DA_FROM</type>
<position>132,99.5</position>
<input>
<ID>IN_0</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>186</ID>
<type>DA_FROM</type>
<position>49.5,-10</position>
<input>
<ID>IN_0</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr4</lparam></gate>
<gate>
<ID>188</ID>
<type>DA_FROM</type>
<position>130.5,64.5</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>189</ID>
<type>DA_FROM</type>
<position>-83,82.5</position>
<input>
<ID>IN_0</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>190</ID>
<type>DA_FROM</type>
<position>130.5,62.5</position>
<input>
<ID>IN_0</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_AND2</type>
<position>135.5,63.5</position>
<input>
<ID>IN_0</ID>117 </input>
<input>
<ID>IN_1</ID>116 </input>
<output>
<ID>OUT</ID>379 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>DA_FROM</type>
<position>46.5,-22</position>
<input>
<ID>IN_0</ID>299 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr15</lparam></gate>
<gate>
<ID>193</ID>
<type>DA_FROM</type>
<position>125.5,57.5</position>
<input>
<ID>IN_0</ID>121 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>346</ID>
<type>DA_FROM</type>
<position>-99.5,99</position>
<input>
<ID>IN_0</ID>224 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>194</ID>
<type>AA_AND3</type>
<position>-72,2.5</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>272 </input>
<input>
<ID>IN_2</ID>352 </input>
<output>
<ID>OUT</ID>340 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>195</ID>
<type>DA_FROM</type>
<position>125.5,55.5</position>
<input>
<ID>IN_0</ID>120 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>356</ID>
<type>DA_FROM</type>
<position>-94.5,92</position>
<input>
<ID>IN_0</ID>243 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>196</ID>
<type>DA_FROM</type>
<position>125.5,52.5</position>
<input>
<ID>IN_0</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>197</ID>
<type>BE_JKFF_LOW</type>
<position>-42,12</position>
<input>
<ID>J</ID>345 </input>
<input>
<ID>K</ID>346 </input>
<output>
<ID>Q</ID>348 </output>
<input>
<ID>clear</ID>351 </input>
<input>
<ID>clock</ID>347 </input>
<output>
<ID>nQ</ID>349 </output>
<input>
<ID>set</ID>351 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>350</ID>
<type>AE_SMALL_INVERTER</type>
<position>-90.5,90</position>
<input>
<ID>IN_0</ID>244 </input>
<output>
<ID>OUT_0</ID>239 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>198</ID>
<type>DA_FROM</type>
<position>125.5,50.5</position>
<input>
<ID>IN_0</ID>118 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>199</ID>
<type>DA_FROM</type>
<position>-22,134</position>
<input>
<ID>IN_0</ID>189 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>344</ID>
<type>AE_OR2</type>
<position>-83.5,101</position>
<input>
<ID>IN_0</ID>226 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>219 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_AND2</type>
<position>130.5,56.5</position>
<input>
<ID>IN_0</ID>121 </input>
<input>
<ID>IN_1</ID>120 </input>
<output>
<ID>OUT</ID>356 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>DA_FROM</type>
<position>-20,127.5</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>354</ID>
<type>AE_SMALL_INVERTER</type>
<position>-90.5,94</position>
<input>
<ID>IN_0</ID>242 </input>
<output>
<ID>OUT_0</ID>241 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>202</ID>
<type>AA_AND2</type>
<position>130.5,51.5</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>118 </input>
<output>
<ID>OUT</ID>355 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>203</ID>
<type>DA_FROM</type>
<position>-81,30.5</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cout</lparam></gate>
<gate>
<ID>364</ID>
<type>FF_GND</type>
<position>88,56</position>
<output>
<ID>OUT_0</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>204</ID>
<type>AE_OR2</type>
<position>139,53.5</position>
<input>
<ID>IN_0</ID>356 </input>
<input>
<ID>IN_1</ID>355 </input>
<output>
<ID>OUT</ID>357 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_AND2</type>
<position>125.5,-47.5</position>
<input>
<ID>IN_0</ID>318 </input>
<input>
<ID>IN_1</ID>319 </input>
<output>
<ID>OUT</ID>322 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>358</ID>
<type>DA_FROM</type>
<position>-94.5,90</position>
<input>
<ID>IN_0</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>206</ID>
<type>DA_FROM</type>
<position>127.5,24.5</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>207</ID>
<type>DA_FROM</type>
<position>-81,-16</position>
<input>
<ID>IN_0</ID>332 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>352</ID>
<type>AA_AND3</type>
<position>-79,88</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>235 </input>
<input>
<ID>IN_2</ID>236 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>208</ID>
<type>DA_FROM</type>
<position>127.5,22.5</position>
<input>
<ID>IN_0</ID>123 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>209</ID>
<type>DA_FROM</type>
<position>24.5,55</position>
<input>
<ID>IN_0</ID>253 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir15</lparam></gate>
<gate>
<ID>362</ID>
<type>AA_AND2</type>
<position>137.5,11</position>
<input>
<ID>IN_0</ID>277 </input>
<input>
<ID>IN_1</ID>282 </input>
<output>
<ID>OUT</ID>279 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_AND2</type>
<position>132.5,23.5</position>
<input>
<ID>IN_0</ID>122 </input>
<input>
<ID>IN_1</ID>123 </input>
<output>
<ID>OUT</ID>314 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>DA_FROM</type>
<position>-22.5,123</position>
<input>
<ID>IN_0</ID>193 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>372</ID>
<type>DA_FROM</type>
<position>53.5,-15.5</position>
<input>
<ID>IN_0</ID>293 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr9</lparam></gate>
<gate>
<ID>212</ID>
<type>AE_OR2</type>
<position>140,25</position>
<input>
<ID>IN_0</ID>313 </input>
<input>
<ID>IN_1</ID>314 </input>
<output>
<ID>OUT</ID>315 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>DA_FROM</type>
<position>-16,101.5</position>
<input>
<ID>IN_0</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID start</lparam></gate>
<gate>
<ID>366</ID>
<type>DA_FROM</type>
<position>120.5,8</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>214</ID>
<type>DA_FROM</type>
<position>120.5,2.5</position>
<input>
<ID>IN_0</ID>128 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>215</ID>
<type>AA_LABEL</type>
<position>62,21.5</position>
<gparam>LABEL_TEXT Check if AC/DR are 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>360</ID>
<type>DA_FROM</type>
<position>-83,80.5</position>
<input>
<ID>IN_0</ID>246 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>216</ID>
<type>DA_FROM</type>
<position>118.5,-56.5</position>
<input>
<ID>IN_0</ID>331 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID start</lparam></gate>
<gate>
<ID>217</ID>
<type>DA_FROM</type>
<position>120.5,-1</position>
<input>
<ID>IN_0</ID>129 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID zeroAC</lparam></gate>
<gate>
<ID>370</ID>
<type>DA_FROM</type>
<position>55.5,-14.5</position>
<input>
<ID>IN_0</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr8</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_AND2</type>
<position>-83.5,108</position>
<input>
<ID>IN_0</ID>220 </input>
<input>
<ID>IN_1</ID>221 </input>
<output>
<ID>OUT</ID>212 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>219</ID>
<type>DA_FROM</type>
<position>120.5,-3</position>
<input>
<ID>IN_0</ID>130 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir2</lparam></gate>
<gate>
<ID>380</ID>
<type>AA_AND2</type>
<position>125.5,-53.5</position>
<input>
<ID>IN_0</ID>327 </input>
<input>
<ID>IN_1</ID>328 </input>
<output>
<ID>OUT</ID>330 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>220</ID>
<type>DA_FROM</type>
<position>-99.5,104</position>
<input>
<ID>IN_0</ID>222 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_AND2</type>
<position>125.5,3.5</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>374</ID>
<type>DA_FROM</type>
<position>120.5,-15</position>
<input>
<ID>IN_0</ID>304 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID zeroDR</lparam></gate>
<gate>
<ID>222</ID>
<type>DA_FROM</type>
<position>-89.5,107</position>
<input>
<ID>IN_0</ID>221 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir7</lparam></gate>
<gate>
<ID>223</ID>
<type>AA_AND2</type>
<position>125.5,-2</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>368</ID>
<type>DE_OR8</type>
<position>62,-9.5</position>
<input>
<ID>IN_0</ID>284 </input>
<input>
<ID>IN_1</ID>285 </input>
<input>
<ID>IN_2</ID>286 </input>
<input>
<ID>IN_3</ID>287 </input>
<input>
<ID>IN_4</ID>291 </input>
<input>
<ID>IN_5</ID>290 </input>
<input>
<ID>IN_6</ID>289 </input>
<input>
<ID>IN_7</ID>288 </input>
<output>
<ID>OUT</ID>283 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>224</ID>
<type>DA_FROM</type>
<position>194.5,119.5</position>
<input>
<ID>IN_0</ID>359 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>225</ID>
<type>DA_FROM</type>
<position>120.5,-8</position>
<input>
<ID>IN_0</ID>133 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir1</lparam></gate>
<gate>
<ID>378</ID>
<type>DA_FROM</type>
<position>120.5,132.5</position>
<input>
<ID>IN_0</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D7</lparam></gate>
<gate>
<ID>226</ID>
<type>DA_FROM</type>
<position>-99.5,102</position>
<input>
<ID>IN_0</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>227</ID>
<type>AA_AND2</type>
<position>125.5,-7</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>260</ID>
<type>DA_FROM</type>
<position>-22,113</position>
<input>
<ID>IN_0</ID>196 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>228</ID>
<type>BE_JKFF_LOW</type>
<position>-67,103</position>
<input>
<ID>J</ID>212 </input>
<input>
<ID>K</ID>219 </input>
<output>
<ID>Q</ID>228 </output>
<input>
<ID>clear</ID>92 </input>
<input>
<ID>clock</ID>210 </input>
<output>
<ID>nQ</ID>229 </output>
<input>
<ID>set</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>229</ID>
<type>AE_OR4</type>
<position>135.5,1.5</position>
<input>
<ID>IN_0</ID>281 </input>
<input>
<ID>IN_1</ID>135 </input>
<input>
<ID>IN_2</ID>137 </input>
<input>
<ID>IN_3</ID>136 </input>
<output>
<ID>OUT</ID>282 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>382</ID>
<type>DA_FROM</type>
<position>118,-54.5</position>
<input>
<ID>IN_0</ID>328 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>230</ID>
<type>DE_TO</type>
<position>214,90.5</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrDR</lparam></gate>
<gate>
<ID>231</ID>
<type>DE_TO</type>
<position>215,109</position>
<input>
<ID>IN_0</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incDR</lparam></gate>
<gate>
<ID>376</ID>
<type>DE_TO</type>
<position>143,-44.5</position>
<input>
<ID>IN_0</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldPC</lparam></gate>
<gate>
<ID>232</ID>
<type>DE_TO</type>
<position>214,97.5</position>
<input>
<ID>IN_0</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID drBus</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_LABEL</type>
<position>23.5,137.5</position>
<gparam>LABEL_TEXT Sequence Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>258</ID>
<type>DA_FROM</type>
<position>-22,130</position>
<input>
<ID>IN_0</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>234</ID>
<type>DA_FROM</type>
<position>194.5,125.5</position>
<input>
<ID>IN_0</ID>363 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>235</ID>
<type>DA_FROM</type>
<position>194.5,121.5</position>
<input>
<ID>IN_0</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>268</ID>
<type>DA_FROM</type>
<position>-5,-21</position>
<input>
<ID>IN_0</ID>375 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir11</lparam></gate>
<gate>
<ID>236</ID>
<type>DA_FROM</type>
<position>194.5,117.5</position>
<input>
<ID>IN_0</ID>361 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>237</ID>
<type>DA_FROM</type>
<position>120.5,-11</position>
<input>
<ID>IN_0</ID>303 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>262</ID>
<type>DA_FROM</type>
<position>-22.5,121</position>
<input>
<ID>IN_0</ID>194 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>238</ID>
<type>DA_FROM</type>
<position>194.5,110</position>
<input>
<ID>IN_0</ID>154 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>239</ID>
<type>AA_AND2</type>
<position>199.5,109</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>155 </input>
<output>
<ID>OUT</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>256</ID>
<type>DA_FROM</type>
<position>-22,132</position>
<input>
<ID>IN_0</ID>191 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>240</ID>
<type>DE_TO</type>
<position>214,-19.5</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrIR</lparam></gate>
<gate>
<ID>241</ID>
<type>DE_TO</type>
<position>213.5,-25.5</position>
<input>
<ID>IN_0</ID>174 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incIR</lparam></gate>
<gate>
<ID>266</ID>
<type>DA_FROM</type>
<position>-5.5,17.5</position>
<input>
<ID>IN_0</ID>208 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>242</ID>
<type>DE_TO</type>
<position>214,-13</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID irBus</lparam></gate>
<gate>
<ID>243</ID>
<type>DA_FROM</type>
<position>198.5,45</position>
<input>
<ID>IN_0</ID>160 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir7</lparam></gate>
<gate>
<ID>276</ID>
<type>DE_TO</type>
<position>5,-7.5</position>
<input>
<ID>IN_0</ID>216 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>244</ID>
<type>AE_OR3</type>
<position>203.5,45</position>
<input>
<ID>IN_0</ID>161 </input>
<input>
<ID>IN_1</ID>160 </input>
<input>
<ID>IN_2</ID>159 </input>
<output>
<ID>OUT</ID>165 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>245</ID>
<type>AA_AND4</type>
<position>211,52</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>1141 </input>
<input>
<ID>IN_2</ID>164 </input>
<input>
<ID>IN_3</ID>165 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>270</ID>
<type>DA_FROM</type>
<position>-8,-2.5</position>
<input>
<ID>IN_0</ID>213 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir9</lparam></gate>
<gate>
<ID>246</ID>
<type>DA_FROM</type>
<position>206,40</position>
<input>
<ID>IN_0</ID>167 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>247</ID>
<type>AA_AND2</type>
<position>211,39</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>166 </input>
<output>
<ID>OUT</ID>170 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>264</ID>
<type>AE_OR2</type>
<position>-17.5,122</position>
<input>
<ID>IN_0</ID>193 </input>
<input>
<ID>IN_1</ID>194 </input>
<output>
<ID>OUT</ID>199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>248</ID>
<type>AE_OR3</type>
<position>220.5,52</position>
<input>
<ID>IN_0</ID>168 </input>
<input>
<ID>IN_1</ID>169 </input>
<input>
<ID>IN_2</ID>170 </input>
<output>
<ID>OUT</ID>1198 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>249</ID>
<type>DA_FROM</type>
<position>210,27</position>
<input>
<ID>IN_0</ID>376 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir5</lparam></gate>
<gate>
<ID>274</ID>
<type>DE_TO</type>
<position>5,-20</position>
<input>
<ID>IN_0</ID>373 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INP</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_AND2</type>
<position>209.5,19.5</position>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>172 </input>
<output>
<ID>OUT</ID>367 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>251</ID>
<type>DA_FROM</type>
<position>204.5,14</position>
<input>
<ID>IN_0</ID>365 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>284</ID>
<type>DE_TO</type>
<position>-59.5,118</position>
<input>
<ID>IN_0</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /FGO</lparam></gate>
<gate>
<ID>252</ID>
<type>DA_FROM</type>
<position>204.5,12</position>
<input>
<ID>IN_0</ID>366 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir10</lparam></gate>
<gate>
<ID>253</ID>
<type>AE_OR2</type>
<position>217,15.5</position>
<input>
<ID>IN_0</ID>367 </input>
<input>
<ID>IN_1</ID>368 </input>
<output>
<ID>OUT</ID>369 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>278</ID>
<type>AA_AND2</type>
<position>0,-1.5</position>
<input>
<ID>IN_0</ID>211 </input>
<input>
<ID>IN_1</ID>213 </input>
<output>
<ID>OUT</ID>214 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>254</ID>
<type>DE_TO</type>
<position>-72,45.5</position>
<input>
<ID>IN_0</ID>323 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrOut</lparam></gate>
<gate>
<ID>255</ID>
<type>DA_FROM</type>
<position>-22,136</position>
<input>
<ID>IN_0</ID>190 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>272</ID>
<type>DE_TO</type>
<position>5,17.5</position>
<input>
<ID>IN_0</ID>208 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>257</ID>
<type>DE_TO</type>
<position>-59,88</position>
<input>
<ID>IN_0</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>259</ID>
<type>DA_FROM</type>
<position>-22.5,117.5</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>261</ID>
<type>AA_AND2</type>
<position>-9,131</position>
<input>
<ID>IN_0</ID>197 </input>
<input>
<ID>IN_1</ID>198 </input>
<output>
<ID>OUT</ID>182 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>263</ID>
<type>AE_OR4</type>
<position>-17,133</position>
<input>
<ID>IN_0</ID>190 </input>
<input>
<ID>IN_1</ID>189 </input>
<input>
<ID>IN_2</ID>191 </input>
<input>
<ID>IN_3</ID>192 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_AND2</type>
<position>-8.5,120.5</position>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_1</ID>200 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>267</ID>
<type>DA_FROM</type>
<position>-13,5</position>
<input>
<ID>IN_0</ID>211 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>269</ID>
<type>DA_FROM</type>
<position>-8,-15</position>
<input>
<ID>IN_0</ID>217 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir6</lparam></gate>
<gate>
<ID>271</ID>
<type>DE_TO</type>
<position>5,22</position>
<input>
<ID>IN_0</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>273</ID>
<type>DE_TO</type>
<position>5,12.5</position>
<input>
<ID>IN_0</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>275</ID>
<type>DE_TO</type>
<position>5,-1.5</position>
<input>
<ID>IN_0</ID>214 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>277</ID>
<type>DE_TO</type>
<position>5,-14</position>
<input>
<ID>IN_0</ID>218 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>279</ID>
<type>AA_AND2</type>
<position>0,-7.5</position>
<input>
<ID>IN_0</ID>211 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>216 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>281</ID>
<type>DA_FROM</type>
<position>-5,-19</position>
<input>
<ID>IN_0</ID>374 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>283</ID>
<type>DA_FROM</type>
<position>121,128.5</position>
<input>
<ID>IN_0</ID>138 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>285</ID>
<type>DA_FROM</type>
<position>-90.5,117</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir10</lparam></gate>
<gate>
<ID>287</ID>
<type>DA_FROM</type>
<position>-74.5,120</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>289</ID>
<type>DE_TO</type>
<position>-58.5,133</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /FGI</lparam></gate>
<gate>
<ID>291</ID>
<type>AA_LABEL</type>
<position>-88.5,140.5</position>
<gparam>LABEL_TEXT fgi</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>AA_LABEL</type>
<position>-88,125</position>
<gparam>LABEL_TEXT fgo</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>295</ID>
<type>DE_TO</type>
<position>-35,10</position>
<input>
<ID>IN_0</ID>349 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /E</lparam></gate>
<gate>
<ID>297</ID>
<type>DE_OR8</type>
<position>62,-18.5</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>293 </input>
<input>
<ID>IN_2</ID>294 </input>
<input>
<ID>IN_3</ID>295 </input>
<input>
<ID>IN_4</ID>299 </input>
<input>
<ID>IN_5</ID>298 </input>
<input>
<ID>IN_6</ID>297 </input>
<input>
<ID>IN_7</ID>296 </input>
<output>
<ID>OUT</ID>300 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>299</ID>
<type>AE_OR2</type>
<position>136.5,-44.5</position>
<input>
<ID>IN_0</ID>321 </input>
<input>
<ID>IN_1</ID>322 </input>
<output>
<ID>OUT</ID>320 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>987</ID>
<type>AA_AND3</type>
<position>125,-20.5</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>306 </input>
<input>
<ID>IN_2</ID>163 </input>
<output>
<ID>OUT</ID>1142 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>301</ID>
<type>DE_TO</type>
<position>-59.5,122</position>
<input>
<ID>IN_0</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGO</lparam></gate>
<gate>
<ID>303</ID>
<type>DA_FROM</type>
<position>-89.5,132</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir11</lparam></gate>
<gate>
<ID>1007</ID>
<type>DA_FROM</type>
<position>-74.5,127</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID start</lparam></gate>
<gate>
<ID>305</ID>
<type>AA_LABEL</type>
<position>-98,148</position>
<gparam>LABEL_TEXT Flags</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>307</ID>
<type>AA_AND3</type>
<position>-6.5,62</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>95 </input>
<input>
<ID>IN_2</ID>96 </input>
<output>
<ID>OUT</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>309</ID>
<type>DA_FROM</type>
<position>-15.5,62</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID I</lparam></gate>
<gate>
<ID>311</ID>
<type>AA_AND3</type>
<position>-6.5,54</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>99 </input>
<input>
<ID>IN_2</ID>100 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>313</ID>
<type>DA_FROM</type>
<position>-15,56</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>315</ID>
<type>DA_FROM</type>
<position>-15,52</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>317</ID>
<type>BE_JKFF_LOW</type>
<position>-67,86</position>
<input>
<ID>J</ID>238 </input>
<input>
<ID>K</ID>248 </input>
<output>
<ID>Q</ID>131 </output>
<input>
<ID>clear</ID>1202 </input>
<input>
<ID>clock</ID>19 </input>
<output>
<ID>nQ</ID>245 </output>
<input>
<ID>set</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>319</ID>
<type>AE_SMALL_INVERTER</type>
<position>-94,6.5</position>
<input>
<ID>IN_0</ID>270 </input>
<output>
<ID>OUT_0</ID>354 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>320</ID>
<type>DA_FROM</type>
<position>49,99.5</position>
<input>
<ID>IN_0</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID start</lparam></gate>
<gate>
<ID>321</ID>
<type>BE_NOR2</type>
<position>75,-15</position>
<input>
<ID>IN_0</ID>283 </input>
<input>
<ID>IN_1</ID>300 </input>
<output>
<ID>OUT</ID>301 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>322</ID>
<type>DA_FROM</type>
<position>50.5,94.5</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir0</lparam></gate>
<gate>
<ID>323</ID>
<type>AE_OR4</type>
<position>199.5,118.5</position>
<input>
<ID>IN_0</ID>360 </input>
<input>
<ID>IN_1</ID>359 </input>
<input>
<ID>IN_2</ID>361 </input>
<input>
<ID>IN_3</ID>358 </input>
<output>
<ID>OUT</ID>362 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>324</ID>
<type>DE_TO</type>
<position>79.5,95.5</position>
<input>
<ID>IN_0</ID>178 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /s</lparam></gate>
<gate>
<ID>325</ID>
<type>DA_FROM</type>
<position>118,-41</position>
<input>
<ID>IN_0</ID>316 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>326</ID>
<type>DA_FROM</type>
<position>63.5,97.5</position>
<input>
<ID>IN_0</ID>173 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>327</ID>
<type>DA_FROM</type>
<position>42.5,52.5</position>
<input>
<ID>IN_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>328</ID>
<type>AA_AND2</type>
<position>56.5,95.5</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>152 </input>
<output>
<ID>OUT</ID>176 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>329</ID>
<type>DA_FROM</type>
<position>-81,-2.5</position>
<input>
<ID>IN_0</ID>273 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>330</ID>
<type>DA_FROM</type>
<position>50.5,96.5</position>
<input>
<ID>IN_0</ID>142 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>331</ID>
<type>DA_FROM</type>
<position>-75,103</position>
<input>
<ID>IN_0</ID>210 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>332</ID>
<type>DE_TO</type>
<position>78,99.5</position>
<input>
<ID>IN_0</ID>177 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s</lparam></gate>
<gate>
<ID>333</ID>
<type>DA_FROM</type>
<position>-99.5,97</position>
<input>
<ID>IN_0</ID>225 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir6</lparam></gate>
<gate>
<ID>335</ID>
<type>DA_FROM</type>
<position>195,96.5</position>
<input>
<ID>IN_0</ID>184 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>336</ID>
<type>DA_FROM</type>
<position>118,-52.5</position>
<input>
<ID>IN_0</ID>327 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>337</ID>
<type>DA_FROM</type>
<position>195,98.5</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>338</ID>
<type>AA_AND2</type>
<position>200,97.5</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>184 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>339</ID>
<type>AA_LABEL</type>
<position>85.5,73.5</position>
<gparam>LABEL_TEXT TR Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>340</ID>
<type>DA_FROM</type>
<position>78,52.5</position>
<input>
<ID>IN_0</ID>234 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>341</ID>
<type>DA_FROM</type>
<position>-89.5,109</position>
<input>
<ID>IN_0</ID>220 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>342</ID>
<type>DE_TO</type>
<position>92,64</position>
<input>
<ID>IN_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldTR</lparam></gate>
<gate>
<ID>343</ID>
<type>DE_TO</type>
<position>-60,105</position>
<input>
<ID>IN_0</ID>228 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IEN</lparam></gate>
<gate>
<ID>345</ID>
<type>AA_AND2</type>
<position>-93.5,103</position>
<input>
<ID>IN_0</ID>222 </input>
<input>
<ID>IN_1</ID>223 </input>
<output>
<ID>OUT</ID>226 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>347</ID>
<type>DA_FROM</type>
<position>-100.5,87</position>
<input>
<ID>IN_0</ID>230 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGI</lparam></gate>
<gate>
<ID>348</ID>
<type>DA_FROM</type>
<position>122,138</position>
<input>
<ID>IN_0</ID>114 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>349</ID>
<type>DA_FROM</type>
<position>-88.5,88</position>
<input>
<ID>IN_0</ID>235 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IEN</lparam></gate>
<gate>
<ID>351</ID>
<type>AA_AND3</type>
<position>-85.5,92</position>
<input>
<ID>IN_0</ID>241 </input>
<input>
<ID>IN_1</ID>240 </input>
<input>
<ID>IN_2</ID>239 </input>
<output>
<ID>OUT</ID>237 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>353</ID>
<type>AE_SMALL_INVERTER</type>
<position>-90.5,92</position>
<input>
<ID>IN_0</ID>243 </input>
<output>
<ID>OUT_0</ID>240 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>355</ID>
<type>DA_FROM</type>
<position>-94.5,94</position>
<input>
<ID>IN_0</ID>242 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>357</ID>
<type>AA_AND2</type>
<position>200.5,-13</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>157 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>359</ID>
<type>AA_AND2</type>
<position>200.5,-5.5</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>148 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>AA_AND2</type>
<position>127.5,17.5</position>
<input>
<ID>IN_0</ID>274 </input>
<input>
<ID>IN_1</ID>275 </input>
<output>
<ID>OUT</ID>276 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>363</ID>
<type>AA_AND2</type>
<position>129.5,9</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>280 </input>
<output>
<ID>OUT</ID>281 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>365</ID>
<type>AE_SMALL_INVERTER</type>
<position>124.5,8</position>
<input>
<ID>IN_0</ID>124 </input>
<output>
<ID>OUT_0</ID>280 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>367</ID>
<type>DA_FROM</type>
<position>55.5,-6</position>
<input>
<ID>IN_0</ID>284 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr0</lparam></gate>
<gate>
<ID>369</ID>
<type>DA_FROM</type>
<position>51,-9</position>
<input>
<ID>IN_0</ID>287 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr3</lparam></gate>
<gate>
<ID>371</ID>
<type>DA_FROM</type>
<position>-16,105.5</position>
<input>
<ID>IN_0</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>373</ID>
<type>DA_FROM</type>
<position>47,-21</position>
<input>
<ID>IN_0</ID>298 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr14</lparam></gate>
<gate>
<ID>375</ID>
<type>DA_FROM</type>
<position>118.5,-46.5</position>
<input>
<ID>IN_0</ID>318 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>377</ID>
<type>AA_AND2</type>
<position>-77,53</position>
<input>
<ID>IN_0</ID>325 </input>
<input>
<ID>IN_1</ID>326 </input>
<output>
<ID>OUT</ID>324 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>379</ID>
<type>AE_OR2</type>
<position>135,-55.5</position>
<input>
<ID>IN_0</ID>330 </input>
<input>
<ID>IN_1</ID>331 </input>
<output>
<ID>OUT</ID>329 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>381</ID>
<type>DA_FROM</type>
<position>132,93.5</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>383</ID>
<type>AA_AND2</type>
<position>137,94.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>384</ID>
<type>DA_FROM</type>
<position>132,95.5</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>386</ID>
<type>DA_FROM</type>
<position>122.5,115</position>
<input>
<ID>IN_0</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>388</ID>
<type>AA_AND3</type>
<position>130.5,130.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>134 </input>
<input>
<ID>IN_2</ID>138 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>390</ID>
<type>AE_OR3</type>
<position>148,130.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>65 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>392</ID>
<type>AA_AND2</type>
<position>134.5,119.5</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>144 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>394</ID>
<type>DA_FROM</type>
<position>115,125</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>396</ID>
<type>DA_FROM</type>
<position>115,121</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>398</ID>
<type>DA_FROM</type>
<position>195.5,-4.5</position>
<input>
<ID>IN_0</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>400</ID>
<type>AE_SMALL_INVERTER</type>
<position>-91,14</position>
<input>
<ID>IN_0</ID>267 </input>
<output>
<ID>OUT_0</ID>353 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>402</ID>
<type>DA_FROM</type>
<position>209,-19.5</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID start</lparam></gate>
<gate>
<ID>404</ID>
<type>DA_FROM</type>
<position>78.5,65</position>
<input>
<ID>IN_0</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_AND2</type>
<position>134.5,43</position>
<input>
<ID>IN_0</ID>380 </input>
<input>
<ID>IN_1</ID>381 </input>
<output>
<ID>OUT</ID>383 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>408</ID>
<type>DE_TO</type>
<position>92,61</position>
<input>
<ID>IN_0</ID>205 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrTR</lparam></gate>
<gate>
<ID>410</ID>
<type>DE_TO</type>
<position>90,51.5</position>
<input>
<ID>IN_0</ID>233 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID trBus</lparam></gate>
<gate>
<ID>412</ID>
<type>DA_FROM</type>
<position>78,50.5</position>
<input>
<ID>IN_0</ID>250 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>414</ID>
<type>DA_FROM</type>
<position>120,-30.5</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>416</ID>
<type>DA_FROM</type>
<position>-16,103.5</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>418</ID>
<type>BE_JKFF_LOW</type>
<position>47.5,58</position>
<input>
<ID>J</ID>254 </input>
<input>
<ID>K</ID>255 </input>
<output>
<ID>Q</ID>257 </output>
<input>
<ID>clear</ID>350 </input>
<input>
<ID>clock</ID>256 </input>
<output>
<ID>nQ</ID>258 </output>
<input>
<ID>set</ID>350 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>419</ID>
<type>AA_AND3</type>
<position>-72,18</position>
<input>
<ID>IN_0</ID>265 </input>
<input>
<ID>IN_1</ID>266 </input>
<input>
<ID>IN_2</ID>267 </input>
<output>
<ID>OUT</ID>338 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>420</ID>
<type>AA_AND3</type>
<position>-72,25</position>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>263 </input>
<input>
<ID>IN_2</ID>264 </input>
<output>
<ID>OUT</ID>337 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>422</ID>
<type>DA_FROM</type>
<position>-81,20</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>424</ID>
<type>DA_FROM</type>
<position>-81,13</position>
<input>
<ID>IN_0</ID>268 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>425</ID>
<type>AA_AND3</type>
<position>-72,-11.5</position>
<input>
<ID>IN_0</ID>310 </input>
<input>
<ID>IN_1</ID>311 </input>
<input>
<ID>IN_2</ID>353 </input>
<output>
<ID>OUT</ID>342 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>426</ID>
<type>DA_FROM</type>
<position>-81,-25</position>
<input>
<ID>IN_0</ID>335 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir10</lparam></gate>
<gate>
<ID>427</ID>
<type>DA_FROM</type>
<position>-81,-4.5</position>
<input>
<ID>IN_0</ID>278 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir8</lparam></gate>
<gate>
<ID>428</ID>
<type>AA_AND2</type>
<position>39,60</position>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>253 </input>
<output>
<ID>OUT</ID>254 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>429</ID>
<type>DA_FROM</type>
<position>23,62.5</position>
<input>
<ID>IN_0</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>430</ID>
<type>AA_INVERTER</type>
<position>30.5,55</position>
<input>
<ID>IN_0</ID>253 </input>
<output>
<ID>OUT_0</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>431</ID>
<type>DE_TO</type>
<position>53.5,60</position>
<input>
<ID>IN_0</ID>257 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID I</lparam></gate>
<gate>
<ID>432</ID>
<type>DA_FROM</type>
<position>-81,23</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /E</lparam></gate>
<gate>
<ID>433</ID>
<type>DA_FROM</type>
<position>-81,-6.5</position>
<input>
<ID>IN_0</ID>309 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>434</ID>
<type>DA_FROM</type>
<position>-81,-22.5</position>
<input>
<ID>IN_0</ID>334 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>435</ID>
<type>DA_FROM</type>
<position>-81,25</position>
<input>
<ID>IN_0</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir8</lparam></gate>
<gate>
<ID>436</ID>
<type>AA_AND3</type>
<position>-72,32.5</position>
<input>
<ID>IN_0</ID>259 </input>
<input>
<ID>IN_1</ID>260 </input>
<input>
<ID>IN_2</ID>261 </input>
<output>
<ID>OUT</ID>336 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>437</ID>
<type>DA_FROM</type>
<position>-81,16</position>
<input>
<ID>IN_0</ID>267 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>438</ID>
<type>DA_FROM</type>
<position>-81,34.5</position>
<input>
<ID>IN_0</ID>259 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>439</ID>
<type>DE_OR8</type>
<position>-56,-3.5</position>
<input>
<ID>IN_0</ID>340 </input>
<input>
<ID>IN_1</ID>341 </input>
<input>
<ID>IN_2</ID>342 </input>
<input>
<ID>IN_3</ID>342 </input>
<input>
<ID>IN_4</ID>987 </input>
<input>
<ID>IN_5</ID>344 </input>
<input>
<ID>IN_6</ID>344 </input>
<input>
<ID>IN_7</ID>343 </input>
<output>
<ID>OUT</ID>346 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>440</ID>
<type>AA_AND3</type>
<position>-72,-18</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>333 </input>
<input>
<ID>IN_2</ID>354 </input>
<output>
<ID>OUT</ID>343 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>441</ID>
<type>DA_FROM</type>
<position>-81,2.5</position>
<input>
<ID>IN_0</ID>272 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>442</ID>
<type>DA_FROM</type>
<position>23,60.5</position>
<input>
<ID>IN_0</ID>251 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>443</ID>
<type>DA_FROM</type>
<position>-81,27</position>
<input>
<ID>IN_0</ID>262 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>444</ID>
<type>DA_FROM</type>
<position>-81,18</position>
<input>
<ID>IN_0</ID>266 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir7</lparam></gate>
<gate>
<ID>445</ID>
<type>AA_AND3</type>
<position>-72,-4.5</position>
<input>
<ID>IN_0</ID>273 </input>
<input>
<ID>IN_1</ID>278 </input>
<input>
<ID>IN_2</ID>309 </input>
<output>
<ID>OUT</ID>341 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>446</ID>
<type>DA_FROM</type>
<position>-81,-9.5</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>447</ID>
<type>DE_TO</type>
<position>-35,14</position>
<input>
<ID>IN_0</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>448</ID>
<type>EE_VDD</type>
<position>47.5,66</position>
<output>
<ID>OUT_0</ID>350 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>450</ID>
<type>AA_AND2</type>
<position>209.5,13</position>
<input>
<ID>IN_0</ID>365 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>368 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>452</ID>
<type>AA_AND2</type>
<position>0,-20</position>
<input>
<ID>IN_0</ID>374 </input>
<input>
<ID>IN_1</ID>375 </input>
<output>
<ID>OUT</ID>373 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>454</ID>
<type>DA_FROM</type>
<position>125.5,44</position>
<input>
<ID>IN_0</ID>380 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>456</ID>
<type>DA_FROM</type>
<position>135.5,38.5</position>
<input>
<ID>IN_0</ID>384 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID start</lparam></gate>
<gate>
<ID>458</ID>
<type>DA_FROM</type>
<position>123,73</position>
<input>
<ID>IN_0</ID>396 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>460</ID>
<type>AE_OR3</type>
<position>144.5,76</position>
<input>
<ID>IN_0</ID>392 </input>
<input>
<ID>IN_1</ID>393 </input>
<input>
<ID>IN_2</ID>394 </input>
<output>
<ID>OUT</ID>391 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>462</ID>
<type>DA_FROM</type>
<position>127,69</position>
<input>
<ID>IN_0</ID>390 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>993</ID>
<type>DA_FROM</type>
<position>206,53</position>
<input>
<ID>IN_0</ID>1141 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /I</lparam></gate>
<gate>
<ID>998</ID>
<type>DA_FROM</type>
<position>120,-26.5</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir8</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_AND3</type>
<position>125,-26.5</position>
<input>
<ID>IN_0</ID>163 </input>
<input>
<ID>IN_1</ID>307 </input>
<input>
<ID>IN_2</ID>104 </input>
<output>
<ID>OUT</ID>308 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_SMALL_INVERTER</type>
<position>-70.5,127</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>1202 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>-72.5,86</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>29</ID>
<type>DA_FROM</type>
<position>-15,97</position>
<input>
<ID>IN_0</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_AND2</type>
<position>-10,96</position>
<input>
<ID>IN_0</ID>249 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>372 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>989</ID>
<type>AE_OR2</type>
<position>2.5,97</position>
<input>
<ID>IN_0</ID>1193 </input>
<input>
<ID>IN_1</ID>372 </input>
<output>
<ID>OUT</ID>1194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>EE_VDD</type>
<position>70.5,103</position>
<output>
<ID>OUT_0</ID>181 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>27 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,121.5,47.5,121.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<connection>
<GID>41</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>155 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,108,196.5,108</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<connection>
<GID>239</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>316 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-41,122.5,-41</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<connection>
<GID>9</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>389 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>129,71,132.5,71</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<connection>
<GID>111</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>30 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,71.5,31.5,71.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<connection>
<GID>63</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>22 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,116.5,58.5,116.5</points>
<connection>
<GID>41</GID>
<name>OUT_1</name></connection>
<connection>
<GID>39</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>317 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-43,122.5,-43</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<connection>
<GID>9</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>385 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>129.5,81.5,132.5,81.5</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<connection>
<GID>459</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,121.5,48.5,124</points>
<connection>
<GID>41</GID>
<name>count_enable</name></connection>
<intersection>124 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,124,48.5,124</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1142 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-24.5,129,-20.5</points>
<intersection>-24.5 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,-20.5,129,-20.5</points>
<connection>
<GID>987</GID>
<name>OUT</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>129,-24.5,130.5,-24.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>129 0</intersection></hsegment></shape></wire>
<wire>
<ID>321 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-43.5,131,-42</points>
<intersection>-43.5 3</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>128.5,-42,131,-42</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131,-43.5,133.5,-43.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>29 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,78.5,31.5,78.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<connection>
<GID>63</GID>
<name>ENABLE</name></connection></hsegment></shape></wire>
<wire>
<ID>23 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,118.5,58.5,118.5</points>
<connection>
<GID>41</GID>
<name>OUT_3</name></connection>
<connection>
<GID>39</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>151 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,101.5,-14,101.5</points>
<connection>
<GID>180</GID>
<name>IN_2</name></connection>
<connection>
<GID>213</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>296 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-19,59,-19</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<connection>
<GID>297</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>351 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42,8,-42,17.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>197</GID>
<name>clear</name></connection>
<connection>
<GID>197</GID>
<name>set</name></connection></vsegment></shape></wire>
<wire>
<ID>32 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,73.5,25.5,74</points>
<intersection>73.5 1</intersection>
<intersection>74 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,73.5,31.5,73.5</points>
<connection>
<GID>63</GID>
<name>IN_2</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,74,25.5,74</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,109,49.5,112.5</points>
<connection>
<GID>41</GID>
<name>clear</name></connection>
<intersection>109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,109,49.5,109</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>315 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,25,143,25</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<connection>
<GID>212</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>163 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120.5,-24.5,120.5,-22.5</points>
<intersection>-24.5 3</intersection>
<intersection>-23.5 4</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120.5,-22.5,122,-22.5</points>
<connection>
<GID>987</GID>
<name>IN_2</name></connection>
<intersection>120.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>120.5,-24.5,122,-24.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>120.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>120,-23.5,120.5,-23.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>120.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>204 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,55,36,55</points>
<connection>
<GID>430</GID>
<name>OUT_0</name></connection>
<connection>
<GID>26</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>12 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,130.5,58.5,130.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>39</GID>
<name>ENABLE</name></connection></hsegment></shape></wire>
<wire>
<ID>333 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,-18,-75,-18</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<connection>
<GID>440</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>269 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,11,-75,11</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<connection>
<GID>391</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>38 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,82,44,82</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>288 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-10,59,-10</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<connection>
<GID>368</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>143 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>117,119,121.5,119</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<connection>
<GID>118</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>15 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,118.5,75.5,118.5</points>
<connection>
<GID>39</GID>
<name>OUT_3</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>235 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-86.5,88,-82,88</points>
<connection>
<GID>352</GID>
<name>IN_1</name></connection>
<connection>
<GID>349</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>268 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,13,-75,13</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<connection>
<GID>424</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>245 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,84,-61,84</points>
<connection>
<GID>317</GID>
<name>nQ</name></connection>
<connection>
<GID>183</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>270 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-94,9,-75,9</points>
<connection>
<GID>15</GID>
<name>IN_2</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-94 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-94,8.5,-94,9</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>9 1</intersection></vsegment></shape></wire>
<wire>
<ID>339 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62.5,11,-62.5,20.5</points>
<intersection>11 2</intersection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62.5,20.5,-59,20.5</points>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<intersection>-62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69,11,-62.5,11</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>-62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-2,130,0.5</points>
<intersection>-2 2</intersection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,0.5,132.5,0.5</points>
<connection>
<GID>229</GID>
<name>IN_2</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128.5,-2,130,-2</points>
<connection>
<GID>223</GID>
<name>OUT</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>290 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,-12,59,-12</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<connection>
<GID>368</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>9 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,122.5,75,122.5</points>
<connection>
<GID>39</GID>
<name>OUT_7</name></connection>
<connection>
<GID>16</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>285 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,-7,59,-7</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<connection>
<GID>368</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>8 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,123.5,80,123.5</points>
<connection>
<GID>39</GID>
<name>OUT_8</name></connection>
<connection>
<GID>54</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>311 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,-11.5,-75,-11.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<connection>
<GID>425</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1198 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223.5,52,223.5,52</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<connection>
<GID>248</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>18 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,115.5,79.5,115.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,127.5,79.5,127.5</points>
<connection>
<GID>39</GID>
<name>OUT_12</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>196 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,113,-20,113</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<connection>
<GID>260</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>3 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>64.5,128.5,75,128.5</points>
<connection>
<GID>39</GID>
<name>OUT_13</name></connection>
<connection>
<GID>49</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>356 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,54.5,135,56.5</points>
<intersection>54.5 2</intersection>
<intersection>56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133.5,56.5,135,56.5</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135,54.5,136,54.5</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>195 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,111,-20,111</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<connection>
<GID>34</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>364 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>211.5,121.5,213.5,121.5</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<connection>
<GID>141</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>203 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,112,-5.5,114.5</points>
<intersection>112 2</intersection>
<intersection>114.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5.5,114.5,5,114.5</points>
<connection>
<GID>42</GID>
<name>IN_2</name></connection>
<intersection>-5.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-14,112,-5.5,112</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,130.5,75,130.5</points>
<connection>
<GID>39</GID>
<name>OUT_15</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>252 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,57,33,61.5</points>
<intersection>57 4</intersection>
<intersection>61 1</intersection>
<intersection>61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,61,36,61</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,61.5,33,61.5</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>33,57,36,57</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>60 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,102.5,141,107</points>
<intersection>102.5 2</intersection>
<intersection>107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,107,141,107</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141,102.5,141.5,102.5</points>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>295 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-17.5,59,-17.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>59 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>59,-18,59,-17.5</points>
<connection>
<GID>297</GID>
<name>IN_3</name></connection>
<intersection>-17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>56 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>140,100.5,141.5,100.5</points>
<connection>
<GID>182</GID>
<name>OUT</name></connection>
<connection>
<GID>385</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>61 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,94.5,141,98.5</points>
<intersection>94.5 1</intersection>
<intersection>98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,94.5,141,94.5</points>
<connection>
<GID>383</GID>
<name>OUT</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141,98.5,141.5,98.5</points>
<connection>
<GID>385</GID>
<name>IN_2</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>272 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,2.5,-75,2.5</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<connection>
<GID>441</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>255 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>42,56,44.5,56</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<connection>
<GID>418</GID>
<name>K</name></connection></hsegment></shape></wire>
<wire>
<ID>63 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147.5,100.5,149.5,100.5</points>
<connection>
<GID>385</GID>
<name>OUT</name></connection>
<connection>
<GID>135</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,117.5,79.5,117.5</points>
<connection>
<GID>39</GID>
<name>OUT_2</name></connection>
<connection>
<GID>60</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>319 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120.5,-48.5,122.5,-48.5</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>233 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,51.5,88,51.5</points>
<connection>
<GID>411</GID>
<name>OUT</name></connection>
<connection>
<GID>410</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>258 </ID>
<shape>
<hsegment>
<ID>10</ID>
<points>50.5,56,51.5,56</points>
<connection>
<GID>418</GID>
<name>nQ</name></connection>
<connection>
<GID>389</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>25 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,112,47.5,112.5</points>
<connection>
<GID>41</GID>
<name>clock</name></connection>
<intersection>112 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,112,47.5,112</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>306 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-20.5,122,-20.5</points>
<connection>
<GID>996</GID>
<name>IN_0</name></connection>
<connection>
<GID>987</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>153 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197.5,-12,197.5,-12</points>
<connection>
<GID>399</GID>
<name>IN_0</name></connection>
<connection>
<GID>357</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>7 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,124.5,75,124.5</points>
<connection>
<GID>39</GID>
<name>OUT_9</name></connection>
<connection>
<GID>33</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>115 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124.5,136,128.5,136</points>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<connection>
<GID>387</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>20 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,95,-13,95</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>50 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,132.5,135,137</points>
<intersection>132.5 1</intersection>
<intersection>137 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,132.5,145,132.5</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>134.5,137,135,137</points>
<connection>
<GID>387</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>114 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,138,128.5,138</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<connection>
<GID>387</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,116.5,76,116.5</points>
<connection>
<GID>39</GID>
<name>OUT_1</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>391 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147.5,76,149,76</points>
<connection>
<GID>460</GID>
<name>OUT</name></connection>
<connection>
<GID>103</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>24 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,115.5,58.5,115.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>21 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,117.5,58.5,117.5</points>
<connection>
<GID>41</GID>
<name>OUT_2</name></connection>
<connection>
<GID>39</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>987 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59,-27.5,-59,-7</points>
<connection>
<GID>439</GID>
<name>IN_4</name></connection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-75.5,-27.5,-59,-27.5</points>
<connection>
<GID>988</GID>
<name>IN_0</name></connection>
<intersection>-59 0</intersection></hsegment></shape></wire>
<wire>
<ID>301 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>78,-15,78.5,-15</points>
<connection>
<GID>321</GID>
<name>OUT</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,125.5,80,125.5</points>
<connection>
<GID>39</GID>
<name>OUT_10</name></connection>
<connection>
<GID>52</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>64.5,126.5,75,126.5</points>
<connection>
<GID>39</GID>
<name>OUT_11</name></connection>
<connection>
<GID>50</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,129.5,79.5,129.5</points>
<connection>
<GID>39</GID>
<name>OUT_14</name></connection>
<connection>
<GID>47</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,119.5,80,119.5</points>
<connection>
<GID>39</GID>
<name>OUT_4</name></connection>
<connection>
<GID>59</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>358 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,115.5,196.5,115.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<connection>
<GID>323</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>205 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>77,61,90,61</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<connection>
<GID>408</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>64.5,120.5,75,120.5</points>
<connection>
<GID>39</GID>
<name>OUT_5</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,121.5,80,121.5</points>
<connection>
<GID>39</GID>
<name>OUT_6</name></connection>
<connection>
<GID>55</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>174 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>209.5,-25.5,211.5,-25.5</points>
<connection>
<GID>401</GID>
<name>OUT_0</name></connection>
<connection>
<GID>241</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>182 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,118.5,-0.5,131</points>
<intersection>118.5 2</intersection>
<intersection>131 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,131,-0.5,131</points>
<connection>
<GID>261</GID>
<name>OUT</name></connection>
<intersection>-0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-0.5,118.5,5,118.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>202 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,116.5,-1.5,120.5</points>
<intersection>116.5 2</intersection>
<intersection>120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5.5,120.5,-1.5,120.5</points>
<connection>
<GID>265</GID>
<name>OUT</name></connection>
<intersection>-1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,116.5,5,116.5</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>-1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>198 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,127.5,-15,130</points>
<intersection>127.5 1</intersection>
<intersection>130 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-18,127.5,-15,127.5</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>-15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15,130,-12,130</points>
<connection>
<GID>261</GID>
<name>IN_1</name></connection>
<intersection>-15 0</intersection></hsegment></shape></wire>
<wire>
<ID>1194 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,97,5,112.5</points>
<connection>
<GID>42</GID>
<name>IN_3</name></connection>
<intersection>97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,97,5.5,97</points>
<connection>
<GID>989</GID>
<name>OUT</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>180 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,115.5,12,115.5</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<connection>
<GID>136</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>140 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>117,123,121.5,123</points>
<connection>
<GID>395</GID>
<name>IN_0</name></connection>
<connection>
<GID>118</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>323 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80,45.5,-74,45.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<connection>
<GID>254</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>188 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81,63,82,63</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<connection>
<GID>403</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1202 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65.5,82,-65.5,131</points>
<intersection>82 9</intersection>
<intersection>116 5</intersection>
<intersection>127 7</intersection>
<intersection>131 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-67,116,-65.5,116</points>
<connection>
<GID>298</GID>
<name>clear</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-67,131,-65.5,131</points>
<connection>
<GID>294</GID>
<name>clear</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-68.5,127,-65.5,127</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-67,82,-65.5,82</points>
<connection>
<GID>317</GID>
<name>clear</name></connection>
<intersection>-65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>206 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,62.5,26.5,62.5</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>284 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-6,59,-6</points>
<connection>
<GID>367</GID>
<name>IN_0</name></connection>
<connection>
<GID>368</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>251 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,60.5,26.5,60.5</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<connection>
<GID>46</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>101 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-32.5,122,-32.5</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<connection>
<GID>413</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>303 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-11,122.5,-11</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<connection>
<GID>237</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>149 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197.5,-4.5,197.5,-4.5</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<connection>
<GID>398</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>302 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-13,122.5,-13</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<connection>
<GID>100</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>159 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200.5,43,200.5,43</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<connection>
<GID>244</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>304 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-15,122.5,-15</points>
<connection>
<GID>48</GID>
<name>IN_2</name></connection>
<connection>
<GID>374</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>305 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-13,145,9</points>
<intersection>-13 2</intersection>
<intersection>9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,9,147,9</points>
<connection>
<GID>119</GID>
<name>IN_2</name></connection>
<intersection>145 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128.5,-13,145,-13</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>145 0</intersection></hsegment></shape></wire>
<wire>
<ID>232 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,57,90,57</points>
<connection>
<GID>364</GID>
<name>OUT_0</name></connection>
<connection>
<GID>409</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>104 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-28.5,122,-28.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<connection>
<GID>123</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>187 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>80.5,65,82,65</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<connection>
<GID>404</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>354 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-94,-20,-94,4.5</points>
<connection>
<GID>319</GID>
<name>OUT_0</name></connection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-94,-20,-75,-20</points>
<connection>
<GID>440</GID>
<name>IN_2</name></connection>
<intersection>-94 0</intersection></hsegment></shape></wire>
<wire>
<ID>201 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,64,90,64</points>
<connection>
<GID>403</GID>
<name>OUT</name></connection>
<connection>
<GID>342</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>249 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,97,-13,97</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>274 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>122,18.5,124.5,18.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<connection>
<GID>361</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>89 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-30.5,122,-30.5</points>
<connection>
<GID>413</GID>
<name>IN_0</name></connection>
<connection>
<GID>414</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>103 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-31.5,129.5,-28.5</points>
<intersection>-31.5 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,-31.5,129.5,-31.5</points>
<connection>
<GID>413</GID>
<name>OUT</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>129.5,-28.5,130.5,-28.5</points>
<connection>
<GID>142</GID>
<name>IN_2</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>334 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,-22.5,-75,-22.5</points>
<connection>
<GID>423</GID>
<name>IN_0</name></connection>
<connection>
<GID>434</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>335 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77,-25,-77,-24.5</points>
<intersection>-25 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-77,-24.5,-75,-24.5</points>
<connection>
<GID>423</GID>
<name>IN_1</name></connection>
<intersection>-77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79,-25,-77,-25</points>
<connection>
<GID>426</GID>
<name>IN_0</name></connection>
<intersection>-77 0</intersection></hsegment></shape></wire>
<wire>
<ID>199 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,121.5,-13,122</points>
<intersection>121.5 1</intersection>
<intersection>122 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,121.5,-11.5,121.5</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-14.5,122,-13,122</points>
<connection>
<GID>264</GID>
<name>OUT</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>344 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60,-23.5,-60,-5</points>
<intersection>-23.5 1</intersection>
<intersection>-6 3</intersection>
<intersection>-5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69,-23.5,-60,-23.5</points>
<connection>
<GID>423</GID>
<name>OUT</name></connection>
<intersection>-60 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-60,-5,-59,-5</points>
<connection>
<GID>439</GID>
<name>IN_6</name></connection>
<intersection>-60 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-60,-6,-59,-6</points>
<connection>
<GID>439</GID>
<name>IN_5</name></connection>
<intersection>-60 0</intersection></hsegment></shape></wire>
<wire>
<ID>352 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88,0.5,-88,24.5</points>
<connection>
<GID>449</GID>
<name>OUT_0</name></connection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-88,0.5,-75,0.5</points>
<connection>
<GID>194</GID>
<name>IN_2</name></connection>
<intersection>-88 0</intersection></hsegment></shape></wire>
<wire>
<ID>207 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3.5,22,3,22</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<connection>
<GID>271</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>347 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-46,12,-45,12</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<connection>
<GID>197</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>329 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>138,-55.5,141,-55.5</points>
<connection>
<GID>379</GID>
<name>OUT</name></connection>
<connection>
<GID>58</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>234 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,52.5,82,52.5</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<connection>
<GID>340</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>250 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,50.5,82,50.5</points>
<connection>
<GID>411</GID>
<name>IN_1</name></connection>
<connection>
<GID>412</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>393 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>138.5,76,141.5,76</points>
<connection>
<GID>306</GID>
<name>OUT</name></connection>
<connection>
<GID>460</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>34 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,78.5,45,78.5</points>
<connection>
<GID>63</GID>
<name>OUT_7</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>37.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37.5,78.5,37.5,82</points>
<intersection>78.5 1</intersection>
<intersection>82 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37.5,82,39,82</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>37.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>271 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,4.5,-75,4.5</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<connection>
<GID>194</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>336 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64,26.5,-64,32.5</points>
<intersection>26.5 1</intersection>
<intersection>32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64,26.5,-59,26.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69,32.5,-64,32.5</points>
<connection>
<GID>436</GID>
<name>OUT</name></connection>
<intersection>-64 0</intersection></hsegment></shape></wire>
<wire>
<ID>337 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64,24.5,-64,25</points>
<intersection>24.5 1</intersection>
<intersection>25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64,24.5,-59,24.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>-64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69,25,-64,25</points>
<connection>
<GID>420</GID>
<name>OUT</name></connection>
<intersection>-64 0</intersection></hsegment></shape></wire>
<wire>
<ID>338 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64,18,-64,22.5</points>
<intersection>18 2</intersection>
<intersection>22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64,22.5,-59,22.5</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<intersection>-64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69,18,-64,18</points>
<connection>
<GID>419</GID>
<name>OUT</name></connection>
<intersection>-64 0</intersection></hsegment></shape></wire>
<wire>
<ID>345 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48.5,14,-48.5,23.5</points>
<intersection>14 1</intersection>
<intersection>23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,14,-45,14</points>
<connection>
<GID>197</GID>
<name>J</name></connection>
<intersection>-48.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52,23.5,-48.5,23.5</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>-48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,72.5,31.5,72.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<connection>
<GID>63</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>33 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,71.5,50.5,71.5</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<connection>
<GID>81</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>41 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,72.5,45,72.5</points>
<connection>
<GID>63</GID>
<name>OUT_1</name></connection>
<connection>
<GID>79</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>40 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,73.5,50.5,73.5</points>
<connection>
<GID>63</GID>
<name>OUT_2</name></connection>
<connection>
<GID>77</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>39 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,74.5,45,74.5</points>
<connection>
<GID>63</GID>
<name>OUT_3</name></connection>
<connection>
<GID>74</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>37 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,75.5,50.5,75.5</points>
<connection>
<GID>63</GID>
<name>OUT_4</name></connection>
<connection>
<GID>72</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>387 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>129,77,132.5,77</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<connection>
<GID>306</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>36 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,76.5,45,76.5</points>
<connection>
<GID>63</GID>
<name>OUT_5</name></connection>
<connection>
<GID>70</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>35 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,77.5,50.5,77.5</points>
<connection>
<GID>63</GID>
<name>OUT_6</name></connection>
<connection>
<GID>68</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>277 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>122.5,12,134.5,12</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>122.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>122.5,12,122.5,12.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>12 1</intersection></vsegment></shape></wire>
<wire>
<ID>275 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>122,16.5,124.5,16.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<connection>
<GID>361</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>377 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212,29,212,29</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<connection>
<GID>453</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>362 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,118.5,204.5,120.5</points>
<intersection>118.5 1</intersection>
<intersection>120.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203.5,118.5,204.5,118.5</points>
<connection>
<GID>323</GID>
<name>OUT</name></connection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>204.5,120.5,205.5,120.5</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>204.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>209 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3.5,12.5,3,12.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<connection>
<GID>273</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>360 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,121.5,196.5,121.5</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<connection>
<GID>323</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>215 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5.5,-8.5,-3,-8.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>325 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80,54,-80,54</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<connection>
<GID>377</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>291 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,-13.5,59,-13.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>59 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>59,-13.5,59,-13</points>
<connection>
<GID>368</GID>
<name>IN_4</name></connection>
<intersection>-13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>313 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,26,135,26.5</points>
<intersection>26 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,26,137,26</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132.5,26.5,135,26.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>167 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,40,208,40</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<connection>
<GID>247</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>312 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154,10,154,10</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<connection>
<GID>119</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>148 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197.5,-6.5,197.5,-6.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<connection>
<GID>359</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>229 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,101,-62,101</points>
<connection>
<GID>228</GID>
<name>nQ</name></connection>
<connection>
<GID>97</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>382 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>146.5,42,147,42</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<connection>
<GID>455</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>150 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>203.5,-5.5,212,-5.5</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<connection>
<GID>359</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>146 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,130.5,154,130.5</points>
<connection>
<GID>390</GID>
<name>OUT</name></connection>
<connection>
<GID>89</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>261 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88,30.5,-75,30.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<connection>
<GID>436</GID>
<name>IN_2</name></connection>
<intersection>-88 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-88,28.5,-88,30.5</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>30.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>395 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131.5,73,132.5,73</points>
<connection>
<GID>463</GID>
<name>OUT_0</name></connection>
<connection>
<GID>111</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>44 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,74.5,207,74.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<connection>
<GID>93</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>45 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,76.5,207,76.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<connection>
<GID>93</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>371 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,74.5,213,75.5</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<intersection>74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213,74.5,213.5,74.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>231 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-98.5,85,-98.5,85</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<connection>
<GID>166</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>376 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212,27,212,27</points>
<connection>
<GID>453</GID>
<name>IN_1</name></connection>
<connection>
<GID>249</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>225 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97.5,97,-96.5,97</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<connection>
<GID>161</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>378 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,28,218,28</points>
<connection>
<GID>453</GID>
<name>OUT</name></connection>
<connection>
<GID>110</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>348 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-39,14,-37,14</points>
<connection>
<GID>197</GID>
<name>Q</name></connection>
<connection>
<GID>447</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1199 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>219.5,73.5,220,73.5</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>396 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,73,127.5,73</points>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<connection>
<GID>463</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>54 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200,67.5,208,67.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>208 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>208,66.5,208,67.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>67.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>92 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68,90,-68,139.5</points>
<intersection>90 2</intersection>
<intersection>99 8</intersection>
<intersection>107 3</intersection>
<intersection>124 5</intersection>
<intersection>139 6</intersection>
<intersection>139.5 7</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-68,90,-67,90</points>
<connection>
<GID>317</GID>
<name>set</name></connection>
<intersection>-68 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-68,107,-67,107</points>
<connection>
<GID>228</GID>
<name>set</name></connection>
<intersection>-68 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-68,124,-67,124</points>
<connection>
<GID>298</GID>
<name>set</name></connection>
<intersection>-68 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-68,139,-67,139</points>
<connection>
<GID>294</GID>
<name>set</name></connection>
<intersection>-68 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-68,139.5,-67,139.5</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<intersection>-68 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-68,99,-67,99</points>
<connection>
<GID>228</GID>
<name>clear</name></connection>
<intersection>-68 0</intersection></hsegment></shape></wire>
<wire>
<ID>217 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,-15,-3,-15</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<connection>
<GID>280</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>370 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213.5,72.5,213.5,72.5</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<connection>
<GID>133</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>93 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3.5,62,0,62</points>
<connection>
<GID>307</GID>
<name>OUT</name></connection>
<connection>
<GID>101</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>386 </ID>
<shape>
<hsegment>
<ID>11</ID>
<points>129.5,79.5,132.5,79.5</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<connection>
<GID>459</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>51 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200.5,65,200.5,65</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<connection>
<GID>108</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>52 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200.5,63,200.5,63</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<connection>
<GID>108</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>388 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>129,75,132.5,75</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<connection>
<GID>306</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>53 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200.5,61,200.5,61</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<connection>
<GID>108</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>392 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,78,140,80.5</points>
<intersection>78 1</intersection>
<intersection>80.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,78,141.5,78</points>
<connection>
<GID>460</GID>
<name>IN_0</name></connection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138.5,80.5,140,80.5</points>
<connection>
<GID>459</GID>
<name>OUT</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>55 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,63,207,64.5</points>
<intersection>63 2</intersection>
<intersection>64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207,64.5,208,64.5</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>206.5,63,207,63</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>168 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215.5,54,215.5,65.5</points>
<intersection>54 3</intersection>
<intersection>65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>214,65.5,215.5,65.5</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<intersection>215.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>215.5,54,217.5,54</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>215.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>390 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>129,69,132.5,69</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<connection>
<GID>111</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>394 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,71,140,74</points>
<intersection>71 2</intersection>
<intersection>74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,74,141.5,74</points>
<connection>
<GID>460</GID>
<name>IN_2</name></connection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138.5,71,140,71</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>164 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,51,208,51</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<connection>
<GID>245</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>314 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,23.5,136.5,24</points>
<intersection>23.5 2</intersection>
<intersection>24 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>135.5,23.5,136.5,23.5</points>
<connection>
<GID>210</GID>
<name>OUT</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>136.5,24,137,24</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200.5,47,200.5,47</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<connection>
<GID>244</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>127 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,4.5,122.5,4.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<connection>
<GID>221</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>126 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>122.5,10,126.5,10</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<connection>
<GID>363</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>132 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-6,122.5,-6</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<connection>
<GID>227</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>300 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-18.5,69,-16</points>
<intersection>-18.5 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-16,72,-16</points>
<connection>
<GID>321</GID>
<name>IN_1</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66,-18.5,69,-18.5</points>
<connection>
<GID>297</GID>
<name>OUT</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>139 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>117,125,121.5,125</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<connection>
<GID>118</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>294 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-16.5,59,-16.5</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>59 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>59,-17,59,-16.5</points>
<connection>
<GID>297</GID>
<name>IN_2</name></connection>
<intersection>-16.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>141 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>117,121,121.5,121</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<connection>
<GID>118</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>106 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,120.5,130,122</points>
<intersection>120.5 1</intersection>
<intersection>122 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,120.5,131.5,120.5</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128.5,122,130,122</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>243 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-92.5,92,-92.5,92</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<connection>
<GID>353</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>276 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,13,141,17.5</points>
<intersection>13 1</intersection>
<intersection>17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141,13,147,13</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>130.5,17.5,141,17.5</points>
<connection>
<GID>361</GID>
<name>OUT</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>279 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>140.5,11,147,11</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<connection>
<GID>362</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>105 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147,-26.5,147,7</points>
<connection>
<GID>119</GID>
<name>IN_3</name></connection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>136.5,-26.5,147,-26.5</points>
<connection>
<GID>142</GID>
<name>OUT</name></connection>
<intersection>147 0</intersection></hsegment></shape></wire>
<wire>
<ID>171 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,20.5,206.5,20.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<connection>
<GID>250</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>369 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,15.5,221.5,15.5</points>
<connection>
<GID>253</GID>
<name>OUT</name></connection>
<connection>
<GID>122</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>172 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,18.5,206.5,18.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<connection>
<GID>250</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>310 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,-9.5,-75,-9.5</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<connection>
<GID>446</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>157 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197.5,-14,197.5,-14</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<connection>
<GID>357</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>166 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,38,208,38</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<connection>
<GID>247</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>227 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88.5,98,-88.5,100</points>
<intersection>98 2</intersection>
<intersection>100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-88.5,100,-86.5,100</points>
<connection>
<GID>344</GID>
<name>IN_1</name></connection>
<intersection>-88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-90.5,98,-88.5,98</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<intersection>-88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>260 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,32.5,-75,32.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<connection>
<GID>436</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>162 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,55,208,55</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<connection>
<GID>245</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>324 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74,53,-74,53</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<connection>
<GID>377</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>46 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-85.5,122,-70,122</points>
<connection>
<GID>292</GID>
<name>OUT_0</name></connection>
<connection>
<GID>298</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>134 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>122.5,130.5,127.5,130.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<connection>
<GID>388</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>42 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-84.5,137,-70,137</points>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection>
<connection>
<GID>294</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>326 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80,52,-80,52</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<connection>
<GID>377</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>372 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7,96,-0.5,96</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<connection>
<GID>989</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>211 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-3,-13,-3,5</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-11,5,-3,5</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>-3 3</intersection></hsegment></shape></wire>
<wire>
<ID>218 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-14,3,-14</points>
<connection>
<GID>280</GID>
<name>OUT</name></connection>
<connection>
<GID>277</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>86 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87.5,134,-86,134</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>379 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>138.5,63.5,141.5,63.5</points>
<connection>
<GID>191</GID>
<name>OUT</name></connection>
<connection>
<GID>137</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>357 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,53.5,144.5,53.5</points>
<connection>
<GID>204</GID>
<name>OUT</name></connection>
<connection>
<GID>138</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>62 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,137,-61,137</points>
<connection>
<GID>294</GID>
<name>Q</name></connection>
<connection>
<GID>300</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>102 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-18.5,122,-18.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<connection>
<GID>987</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>67 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80,133,-70,133</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<connection>
<GID>294</GID>
<name>K</name></connection></hsegment></shape></wire>
<wire>
<ID>49 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-72.5,135,-70,135</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<connection>
<GID>294</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>66 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,133,-60.5,133</points>
<connection>
<GID>294</GID>
<name>nQ</name></connection>
<connection>
<GID>289</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>147 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195.5,90.5,212,90.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<connection>
<GID>230</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>308 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-26.5,130.5,-26.5</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<connection>
<GID>142</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>88 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,119,-87,119</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<connection>
<GID>304</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>363 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,122.5,201,125.5</points>
<intersection>122.5 2</intersection>
<intersection>125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>196.5,125.5,201,125.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>201,122.5,205.5,122.5</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>201 0</intersection></hsegment></shape></wire>
<wire>
<ID>91 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-81,118,-70,118</points>
<connection>
<GID>304</GID>
<name>OUT</name></connection>
<connection>
<GID>298</GID>
<name>K</name></connection></hsegment></shape></wire>
<wire>
<ID>57 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-72.5,120,-70,120</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<connection>
<GID>298</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>59 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,122,-61.5,122</points>
<connection>
<GID>298</GID>
<name>Q</name></connection>
<connection>
<GID>301</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>58 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,118,-61.5,118</points>
<connection>
<GID>298</GID>
<name>nQ</name></connection>
<connection>
<GID>284</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>110 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,108,132.5,109</points>
<intersection>108 2</intersection>
<intersection>109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,109,132.5,109</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132.5,108,134,108</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>111 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,105,132.5,106</points>
<intersection>105 1</intersection>
<intersection>106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,105,132.5,105</points>
<connection>
<GID>179</GID>
<name>OUT</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132.5,106,134,106</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,7.5,59,7.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<connection>
<GID>152</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>94 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,64,-9.5,64</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<connection>
<GID>307</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>383 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137.5,43,140.5,43</points>
<connection>
<GID>406</GID>
<name>OUT</name></connection>
<connection>
<GID>147</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>384 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,38.5,139,41</points>
<intersection>38.5 2</intersection>
<intersection>41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139,41,140.5,41</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137.5,38.5,139,38.5</points>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>76 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,4.5,59,4.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<connection>
<GID>148</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>77 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,3.5,59,3.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<connection>
<GID>148</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>78 </ID>
<shape>
<hsegment>
<ID>9</ID>
<points>54,2.5,59,2.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<connection>
<GID>148</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>79 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,1.5,59,1.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<connection>
<GID>148</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>83 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-2.5,59,-2.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<connection>
<GID>148</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>82 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,-1.5,59,-1.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<connection>
<GID>148</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>81 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-0.5,59,-0.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<connection>
<GID>148</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>80 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,0.5,59,0.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<connection>
<GID>148</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>84 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,1,69,3.5</points>
<intersection>1 2</intersection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,3.5,72,3.5</points>
<connection>
<GID>154</GID>
<name>IN_1</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66,1,69,1</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>87 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87.5,132,-86,132</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>381 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,42,131.5,42</points>
<connection>
<GID>406</GID>
<name>IN_1</name></connection>
<connection>
<GID>149</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>70 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,11.5,59,11.5</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<connection>
<GID>152</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>68 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>57.5,13.5,59,13.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<connection>
<GID>152</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>69 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,12.5,59,12.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<connection>
<GID>152</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>71 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,10.5,59,10.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<connection>
<GID>152</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>75 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,6,59,6</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>59 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>59,6,59,6.5</points>
<connection>
<GID>152</GID>
<name>IN_4</name></connection>
<intersection>6 1</intersection></vsegment></shape></wire>
<wire>
<ID>73 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,8.5,59,8.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<connection>
<GID>152</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>72 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,9.5,59,9.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<connection>
<GID>152</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>43 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,5.5,69,10</points>
<intersection>5.5 1</intersection>
<intersection>10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,5.5,72,5.5</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66,10,69,10</points>
<connection>
<GID>152</GID>
<name>OUT</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>85 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,4.5,79,4.5</points>
<connection>
<GID>154</GID>
<name>OUT</name></connection>
<connection>
<GID>171</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>264 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,23,-75,23</points>
<connection>
<GID>420</GID>
<name>IN_2</name></connection>
<connection>
<GID>432</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>247 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81,82.5,-81,82.5</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<connection>
<GID>189</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>246 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81,80.5,-81,80.5</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<connection>
<GID>360</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>248 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-71.5,81.5,-71.5,84</points>
<intersection>81.5 2</intersection>
<intersection>84 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71.5,84,-70,84</points>
<connection>
<GID>317</GID>
<name>K</name></connection>
<intersection>-71.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-75,81.5,-71.5,81.5</points>
<connection>
<GID>316</GID>
<name>OUT</name></connection>
<intersection>-71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,60,-9.5,60</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<connection>
<GID>307</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>90 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,117,-87,117</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<connection>
<GID>304</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>99 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,54,-9.5,54</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<connection>
<GID>311</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>224 </ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-97.5,99,-96.5,99</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<connection>
<GID>161</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>175 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51,99.5,67.5,99.5</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<connection>
<GID>318</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>176 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,95.5,67.5,95.5</points>
<connection>
<GID>328</GID>
<name>OUT</name></connection>
<connection>
<GID>318</GID>
<name>K</name></connection></hsegment></shape></wire>
<wire>
<ID>181 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,93.5,70.5,102</points>
<connection>
<GID>318</GID>
<name>clear</name></connection>
<connection>
<GID>318</GID>
<name>set</name></connection>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>173 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65.5,97.5,67.5,97.5</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<connection>
<GID>318</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>177 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,99.5,76,99.5</points>
<connection>
<GID>318</GID>
<name>Q</name></connection>
<connection>
<GID>332</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>178 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,95.5,77.5,95.5</points>
<connection>
<GID>318</GID>
<name>nQ</name></connection>
<connection>
<GID>324</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>230 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-98.5,87,-98.5,87</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<connection>
<GID>347</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>236 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-92.5,86,-82,86</points>
<connection>
<GID>166</GID>
<name>OUT</name></connection>
<connection>
<GID>352</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>97 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3.5,54,0.5,54</points>
<connection>
<GID>311</GID>
<name>OUT</name></connection>
<connection>
<GID>312</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>297 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-20,59,-20</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<connection>
<GID>297</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>133 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-8,122.5,-8</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<connection>
<GID>227</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>286 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-8,59,-8</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<connection>
<GID>368</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>108 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,106,125,106</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<connection>
<GID>179</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>109 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,104,125,104</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<connection>
<GID>179</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>107 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,105.5,-14,105.5</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<connection>
<GID>371</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>298 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,-21,59,-21</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<connection>
<GID>297</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>145 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,103.5,-14,103.5</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<connection>
<GID>416</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>350 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,54,47.5,65</points>
<connection>
<GID>448</GID>
<name>OUT_0</name></connection>
<connection>
<GID>418</GID>
<name>set</name></connection>
<connection>
<GID>418</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>197 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,132,-12,133</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>133 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,133,-12,133</points>
<connection>
<GID>263</GID>
<name>OUT</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>1193 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,98,-4,103.5</points>
<intersection>98 1</intersection>
<intersection>103.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,98,-0.5,98</points>
<connection>
<GID>989</GID>
<name>IN_0</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,103.5,-4,103.5</points>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>289 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-11,59,-11</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<connection>
<GID>368</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>112 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,101.5,134,101.5</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<connection>
<GID>184</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>113 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,99.5,134,99.5</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<connection>
<GID>185</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>117 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,64.5,132.5,64.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<connection>
<GID>191</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>116 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,62.5,132.5,62.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<connection>
<GID>191</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>299 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-22,59,-22</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<connection>
<GID>297</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>121 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,57.5,127.5,57.5</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<connection>
<GID>200</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>340 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64,0,-64,2.5</points>
<intersection>0 1</intersection>
<intersection>2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64,0,-59,0</points>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<intersection>-64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69,2.5,-64,2.5</points>
<connection>
<GID>194</GID>
<name>OUT</name></connection>
<intersection>-64 0</intersection></hsegment></shape></wire>
<wire>
<ID>120 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,55.5,127.5,55.5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<connection>
<GID>200</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>119 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,52.5,127.5,52.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<connection>
<GID>202</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>244 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-92.5,90,-92.5,90</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<connection>
<GID>358</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>256 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,52.5,44.5,58</points>
<connection>
<GID>418</GID>
<name>clock</name></connection>
<connection>
<GID>327</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>239 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88.5,90,-88.5,90</points>
<connection>
<GID>350</GID>
<name>OUT_0</name></connection>
<connection>
<GID>351</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>193 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,123,-20.5,123</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<connection>
<GID>264</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>346 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48.5,-3.5,-48.5,10</points>
<intersection>-3.5 2</intersection>
<intersection>10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,10,-45,10</points>
<connection>
<GID>197</GID>
<name>K</name></connection>
<intersection>-48.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52,-3.5,-48.5,-3.5</points>
<connection>
<GID>439</GID>
<name>OUT</name></connection>
<intersection>-48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>349 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-39,10,-37,10</points>
<connection>
<GID>197</GID>
<name>nQ</name></connection>
<connection>
<GID>295</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>118 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,50.5,127.5,50.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<connection>
<GID>202</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>226 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88.5,102,-88.5,103</points>
<intersection>102 1</intersection>
<intersection>103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-88.5,102,-86.5,102</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>-88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-90.5,103,-88.5,103</points>
<connection>
<GID>345</GID>
<name>OUT</name></connection>
<intersection>-88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>380 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,44,131.5,44</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<connection>
<GID>406</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>219 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80.5,101,-70,101</points>
<connection>
<GID>344</GID>
<name>OUT</name></connection>
<connection>
<GID>228</GID>
<name>K</name></connection></hsegment></shape></wire>
<wire>
<ID>189 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,134,-20,134</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<connection>
<GID>263</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>242 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-92.5,94,-92.5,94</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<connection>
<GID>355</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>266 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,18,-75,18</points>
<connection>
<GID>419</GID>
<name>IN_1</name></connection>
<connection>
<GID>444</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>241 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88.5,94,-88.5,94</points>
<connection>
<GID>354</GID>
<name>OUT_0</name></connection>
<connection>
<GID>351</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>355 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,51.5,135,52.5</points>
<intersection>51.5 1</intersection>
<intersection>52.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133.5,51.5,135,51.5</points>
<connection>
<GID>202</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135,52.5,136,52.5</points>
<connection>
<GID>204</GID>
<name>IN_1</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>165 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,45,208,49</points>
<connection>
<GID>245</GID>
<name>IN_3</name></connection>
<intersection>45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>206.5,45,208,45</points>
<connection>
<GID>244</GID>
<name>OUT</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>318 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120.5,-46.5,122.5,-46.5</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<connection>
<GID>205</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>322 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-47.5,131,-45.5</points>
<intersection>-47.5 2</intersection>
<intersection>-45.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>128.5,-47.5,131,-47.5</points>
<connection>
<GID>205</GID>
<name>OUT</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131,-45.5,133.5,-45.5</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>122 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,24.5,129.5,24.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<connection>
<GID>210</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>262 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,27,-75,27</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<connection>
<GID>443</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>237 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-82,90,-82,92</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-82.5,92,-82,92</points>
<connection>
<GID>351</GID>
<name>OUT</name></connection>
<intersection>-82 0</intersection></hsegment></shape></wire>
<wire>
<ID>238 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76,88,-70,88</points>
<connection>
<GID>317</GID>
<name>J</name></connection>
<connection>
<GID>352</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>332 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,-16,-75,-16</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<connection>
<GID>440</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>123 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,22.5,129.5,22.5</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<connection>
<GID>210</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>129 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-1,122.5,-1</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<connection>
<GID>223</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>282 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,1.5,138,10</points>
<intersection>1.5 2</intersection>
<intersection>10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134.5,10,138,10</points>
<connection>
<GID>362</GID>
<name>IN_1</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,1.5,139.5,1.5</points>
<connection>
<GID>229</GID>
<name>OUT</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>278 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,-4.5,-75,-4.5</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<connection>
<GID>445</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>253 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,55,27.5,55</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>27 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>27,55,27,59</points>
<intersection>55 1</intersection>
<intersection>59 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>27,59,36,59</points>
<connection>
<GID>428</GID>
<name>IN_1</name></connection>
<intersection>27 5</intersection></hsegment></shape></wire>
<wire>
<ID>293 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,-15.5,59,-15.5</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>59 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>59,-16,59,-15.5</points>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>-15.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>124 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,8,122.5,8</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<connection>
<GID>365</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>128 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,2.5,122.5,2.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<connection>
<GID>221</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>331 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120.5,-56.5,132,-56.5</points>
<connection>
<GID>379</GID>
<name>IN_1</name></connection>
<connection>
<GID>216</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>131 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,88,-61,88</points>
<connection>
<GID>317</GID>
<name>Q</name></connection>
<connection>
<GID>257</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>292 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-14.5,59,-14.5</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<intersection>59 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>59,-15,59,-14.5</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>220 </ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-87.5,109,-86.5,109</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<connection>
<GID>218</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>374 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-19,-3,-19</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<connection>
<GID>452</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>221 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87.5,107,-86.5,107</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<connection>
<GID>218</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>212 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75.5,105,-75.5,108</points>
<intersection>105 1</intersection>
<intersection>108 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-75.5,105,-70,105</points>
<connection>
<GID>228</GID>
<name>J</name></connection>
<intersection>-75.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-80.5,108,-75.5,108</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<intersection>-75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>327 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>120,-52.5,122.5,-52.5</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<connection>
<GID>380</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>328 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-54.5,122.5,-54.5</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<connection>
<GID>380</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>330 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-54.5,130,-53.5</points>
<intersection>-54.5 1</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-54.5,132,-54.5</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128.5,-53.5,130,-53.5</points>
<connection>
<GID>380</GID>
<name>OUT</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>130 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-3,122.5,-3</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<connection>
<GID>223</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>222 </ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-97.5,104,-96.5,104</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<connection>
<GID>345</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>280 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,8,126.5,8</points>
<connection>
<GID>363</GID>
<name>IN_1</name></connection>
<connection>
<GID>365</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>135 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,2.5,130.5,3.5</points>
<intersection>2.5 1</intersection>
<intersection>3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,2.5,132.5,2.5</points>
<connection>
<GID>229</GID>
<name>IN_1</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128.5,3.5,130.5,3.5</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>287 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-9,59,-9</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<connection>
<GID>368</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>283 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-14,69,-9.5</points>
<intersection>-14 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-14,72,-14</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66,-9.5,69,-9.5</points>
<connection>
<GID>368</GID>
<name>OUT</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>359 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,119.5,196.5,119.5</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<connection>
<GID>323</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>125 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>122.5,132.5,127.5,132.5</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<connection>
<GID>388</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>368 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,13,213,14.5</points>
<intersection>13 1</intersection>
<intersection>14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>212.5,13,213,13</points>
<connection>
<GID>450</GID>
<name>OUT</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213,14.5,214,14.5</points>
<connection>
<GID>253</GID>
<name>IN_1</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>223 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97.5,102,-96.5,102</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<connection>
<GID>345</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>136 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-7,130.5,-1.5</points>
<intersection>-7 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128.5,-7,130.5,-7</points>
<connection>
<GID>227</GID>
<name>OUT</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>130.5,-1.5,132.5,-1.5</points>
<connection>
<GID>229</GID>
<name>IN_3</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>210 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-73,103,-70,103</points>
<connection>
<GID>228</GID>
<name>clock</name></connection>
<connection>
<GID>331</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>228 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,105,-62,105</points>
<connection>
<GID>228</GID>
<name>Q</name></connection>
<connection>
<GID>343</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>281 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,4.5,132.5,9</points>
<connection>
<GID>363</GID>
<name>OUT</name></connection>
<connection>
<GID>229</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>320 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>139.5,-44.5,141,-44.5</points>
<connection>
<GID>299</GID>
<name>OUT</name></connection>
<connection>
<GID>376</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>156 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202.5,109,213,109</points>
<connection>
<GID>239</GID>
<name>OUT</name></connection>
<connection>
<GID>231</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>185 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>203,97.5,212,97.5</points>
<connection>
<GID>338</GID>
<name>OUT</name></connection>
<connection>
<GID>232</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>192 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,130,-20,130</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<connection>
<GID>263</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>375 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-21,-3,-21</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<connection>
<GID>452</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>361 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,117.5,196.5,117.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<connection>
<GID>323</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>194 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,121,-20.5,121</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<connection>
<GID>264</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>154 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,110,196.5,110</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<connection>
<GID>239</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>191 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,132,-20,132</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<connection>
<GID>263</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>186 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>211,-19.5,212,-19.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<connection>
<GID>402</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>208 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3.5,17.5,3,17.5</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<connection>
<GID>272</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>158 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>203.5,-13,212,-13</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<connection>
<GID>357</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>216 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-7.5,3,-7.5</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>160 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200.5,45,200.5,45</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<connection>
<GID>244</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>366 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,12,206.5,12</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<connection>
<GID>450</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>213 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,-2.5,-3,-2.5</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<connection>
<GID>278</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1141 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,53,208,53</points>
<connection>
<GID>245</GID>
<name>IN_1</name></connection>
<connection>
<GID>993</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>169 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>214,52,217.5,52</points>
<connection>
<GID>245</GID>
<name>OUT</name></connection>
<connection>
<GID>248</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>170 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215.5,39,215.5,50</points>
<intersection>39 1</intersection>
<intersection>50 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>214,39,215.5,39</points>
<connection>
<GID>247</GID>
<name>OUT</name></connection>
<intersection>215.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>215.5,50,217.5,50</points>
<connection>
<GID>248</GID>
<name>IN_2</name></connection>
<intersection>215.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>373 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-20,3,-20</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<connection>
<GID>452</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>367 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,16.5,213,19.5</points>
<intersection>16.5 2</intersection>
<intersection>19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>212.5,19.5,213,19.5</points>
<connection>
<GID>250</GID>
<name>OUT</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213,16.5,214,16.5</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>365 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,14,206.5,14</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<connection>
<GID>450</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>214 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-1.5,3,-1.5</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<connection>
<GID>275</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>190 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,136,-20,136</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<connection>
<GID>263</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>200 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,117.5,-16,119.5</points>
<intersection>117.5 1</intersection>
<intersection>119.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20.5,117.5,-16,117.5</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-16,119.5,-11.5,119.5</points>
<connection>
<GID>265</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>138 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,128.5,127.5,128.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<connection>
<GID>388</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>11 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72.5,127,-72.5,127</points>
<connection>
<GID>1007</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>95 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,62,-9.5,62</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<connection>
<GID>307</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>98 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,56,-9.5,56</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<connection>
<GID>311</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>100 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,52,-9.5,52</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<connection>
<GID>311</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>19 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-70.5,86,-70,86</points>
<connection>
<GID>317</GID>
<name>clock</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>152 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,94.5,53.5,94.5</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<connection>
<GID>328</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>142 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,96.5,53.5,96.5</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<connection>
<GID>328</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>273 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,-2.5,-75,-2.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<connection>
<GID>445</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>184 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,96.5,197,96.5</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<connection>
<GID>338</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>183 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,98.5,197,98.5</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<connection>
<GID>338</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>240 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88.5,92,-88.5,92</points>
<connection>
<GID>351</GID>
<name>IN_1</name></connection>
<connection>
<GID>353</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>47 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,93.5,134,93.5</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<connection>
<GID>383</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>48 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,95.5,134,95.5</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<connection>
<GID>384</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>144 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,115,131,118.5</points>
<intersection>115 2</intersection>
<intersection>118.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,118.5,131.5,118.5</points>
<connection>
<GID>392</GID>
<name>IN_1</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,115,131,115</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>64 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,130.5,145,130.5</points>
<connection>
<GID>388</GID>
<name>OUT</name></connection>
<connection>
<GID>390</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>65 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,119.5,139,128.5</points>
<intersection>119.5 5</intersection>
<intersection>128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139,128.5,145,128.5</points>
<connection>
<GID>390</GID>
<name>IN_2</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>137.5,119.5,139,119.5</points>
<connection>
<GID>392</GID>
<name>OUT</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>267 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-91,16,-75,16</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<connection>
<GID>419</GID>
<name>IN_2</name></connection>
<connection>
<GID>437</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>353 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-91,-13.5,-91,12</points>
<connection>
<GID>400</GID>
<name>OUT_0</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-91,-13.5,-75,-13.5</points>
<connection>
<GID>425</GID>
<name>IN_2</name></connection>
<intersection>-91 0</intersection></hsegment></shape></wire>
<wire>
<ID>254 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42,60,44.5,60</points>
<connection>
<GID>428</GID>
<name>OUT</name></connection>
<connection>
<GID>418</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>257 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>50.5,60,51.5,60</points>
<connection>
<GID>418</GID>
<name>Q</name></connection>
<connection>
<GID>431</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>265 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,20,-75,20</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<connection>
<GID>422</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>263 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,25,-75,25</points>
<connection>
<GID>420</GID>
<name>IN_1</name></connection>
<connection>
<GID>435</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>342 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,-11.5,-63.5,-3</points>
<intersection>-11.5 2</intersection>
<intersection>-3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,-3,-59,-3</points>
<connection>
<GID>439</GID>
<name>IN_3</name></connection>
<intersection>-63.5 0</intersection>
<intersection>-59 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69,-11.5,-63.5,-11.5</points>
<connection>
<GID>425</GID>
<name>OUT</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-59,-3,-59,-2</points>
<connection>
<GID>439</GID>
<name>IN_2</name></connection>
<intersection>-3 1</intersection></vsegment></shape></wire>
<wire>
<ID>309 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,-6.5,-75,-6.5</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<connection>
<GID>445</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>259 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,34.5,-75,34.5</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<connection>
<GID>438</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>341 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64,-4.5,-64,-1</points>
<intersection>-4.5 2</intersection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64,-1,-59,-1</points>
<connection>
<GID>439</GID>
<name>IN_1</name></connection>
<intersection>-64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69,-4.5,-64,-4.5</points>
<connection>
<GID>445</GID>
<name>OUT</name></connection>
<intersection>-64 0</intersection></hsegment></shape></wire>
<wire>
<ID>343 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-61.5,-18,-61.5,-4</points>
<intersection>-18 1</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69,-18,-61.5,-18</points>
<connection>
<GID>440</GID>
<name>OUT</name></connection>
<intersection>-61.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-61.5,-4,-59,-4</points>
<connection>
<GID>439</GID>
<name>IN_7</name></connection>
<intersection>-61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>307 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-26.5,122,-26.5</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<connection>
<GID>998</GID>
<name>IN_0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-46.9346,16.0812,95.1634,-53.4409</PageViewport>
<gate>
<ID>513</ID>
<type>DA_FROM</type>
<position>40.5,33.5</position>
<input>
<ID>IN_0</ID>436 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>464</ID>
<type>FF_GND</type>
<position>35.5,26.5</position>
<output>
<ID>OUT_0</ID>445 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>641</ID>
<type>DA_FROM</type>
<position>-65,-38</position>
<input>
<ID>IN_0</ID>686 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>794</ID>
<type>DA_FROM</type>
<position>117,-57</position>
<input>
<ID>IN_0</ID>546 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr11</lparam></gate>
<gate>
<ID>521</ID>
<type>DE_TO</type>
<position>48,-29</position>
<input>
<ID>IN_0</ID>476 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin2</lparam></gate>
<gate>
<ID>472</ID>
<type>DA_FROM</type>
<position>-38.5,-13.5</position>
<input>
<ID>IN_0</ID>418 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>649</ID>
<type>DA_FROM</type>
<position>115.5,18</position>
<input>
<ID>IN_0</ID>559 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum8</lparam></gate>
<gate>
<ID>802</ID>
<type>BV_4x1_BUS_END</type>
<position>-71.5,8.5</position>
<input>
<ID>IN_0</ID>740 </input>
<input>
<ID>IN_1</ID>738 </input>
<input>
<ID>IN_2</ID>739 </input>
<input>
<ID>IN_3</ID>737 </input>
<input>
<ID>OUT</ID>746 747 748 749 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>465</ID>
<type>DA_FROM</type>
<position>-38.5,-21.5</position>
<input>
<ID>IN_0</ID>422 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>631</ID>
<type>AE_SMALL_INVERTER</type>
<position>123.5,0</position>
<input>
<ID>IN_0</ID>577 </input>
<output>
<ID>OUT_0</ID>568 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>466</ID>
<type>DA_FROM</type>
<position>-38.5,-19.5</position>
<input>
<ID>IN_0</ID>421 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>805</ID>
<type>DE_TO</type>
<position>-25,38</position>
<input>
<ID>IN_0</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr15</lparam></gate>
<gate>
<ID>467</ID>
<type>DE_TO</type>
<position>47.5,23</position>
<input>
<ID>IN_0</ID>446 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin0</lparam></gate>
<gate>
<ID>798</ID>
<type>DA_FROM</type>
<position>160.5,-57.5</position>
<input>
<ID>IN_0</ID>606 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr15</lparam></gate>
<gate>
<ID>645</ID>
<type>AE_SMALL_INVERTER</type>
<position>123.5,-28</position>
<input>
<ID>IN_0</ID>592 </input>
<output>
<ID>OUT_0</ID>583 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>468</ID>
<type>DA_FROM</type>
<position>-38.5,-17.5</position>
<input>
<ID>IN_0</ID>420 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INP</lparam></gate>
<gate>
<ID>517</ID>
<type>DA_FROM</type>
<position>24,-8</position>
<input>
<ID>IN_0</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>469</ID>
<type>FF_GND</type>
<position>36,2.5</position>
<output>
<ID>OUT_0</ID>460 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>619</ID>
<type>DA_FROM</type>
<position>93.5,-45.5</position>
<input>
<ID>IN_0</ID>539 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>470</ID>
<type>DA_FROM</type>
<position>-38.5,-15.5</position>
<input>
<ID>IN_0</ID>419 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>793</ID>
<type>DA_FROM</type>
<position>116,-30</position>
<input>
<ID>IN_0</ID>531 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr10</lparam></gate>
<gate>
<ID>471</ID>
<type>DE_TO</type>
<position>48,-1</position>
<input>
<ID>IN_0</ID>461 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin1</lparam></gate>
<gate>
<ID>473</ID>
<type>AI_MUX_8x1</type>
<position>43,-1</position>
<input>
<ID>IN_0</ID>447 </input>
<input>
<ID>IN_1</ID>454 </input>
<input>
<ID>IN_2</ID>455 </input>
<input>
<ID>IN_3</ID>414 </input>
<input>
<ID>IN_4</ID>448 </input>
<input>
<ID>IN_5</ID>458 </input>
<input>
<ID>IN_6</ID>459 </input>
<input>
<ID>IN_7</ID>460 </input>
<output>
<ID>OUT</ID>461 </output>
<input>
<ID>SEL_0</ID>449 </input>
<input>
<ID>SEL_1</ID>450 </input>
<input>
<ID>SEL_2</ID>451 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>639</ID>
<type>AA_AND2</type>
<position>123,14.5</position>
<input>
<ID>IN_0</ID>558 </input>
<input>
<ID>IN_1</ID>557 </input>
<output>
<ID>OUT</ID>552 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>474</ID>
<type>DA_FROM</type>
<position>-38.5,-11.5</position>
<input>
<ID>IN_0</ID>417 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>813</ID>
<type>FF_GND</type>
<position>-39.5,20.5</position>
<output>
<ID>OUT_0</ID>736 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>475</ID>
<type>AE_SMALL_INVERTER</type>
<position>31.5,0</position>
<input>
<ID>IN_0</ID>457 </input>
<output>
<ID>OUT_0</ID>448 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>518</ID>
<type>DA_FROM</type>
<position>45,9.5</position>
<input>
<ID>IN_0</ID>449 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>806</ID>
<type>DE_TO</type>
<position>-25,36</position>
<input>
<ID>IN_0</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr14</lparam></gate>
<gate>
<ID>653</ID>
<type>DE_TO</type>
<position>-8.5,-58</position>
<input>
<ID>IN_0</ID>726 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum0</lparam></gate>
<gate>
<ID>476</ID>
<type>DE_TO</type>
<position>-8.5,-23</position>
<input>
<ID>IN_0</ID>427 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>525</ID>
<type>DA_FROM</type>
<position>24,-36</position>
<input>
<ID>IN_0</ID>468 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>477</ID>
<type>DA_FROM</type>
<position>24,-6</position>
<input>
<ID>IN_0</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum1</lparam></gate>
<gate>
<ID>627</ID>
<type>FF_GND</type>
<position>128,2.5</position>
<output>
<ID>OUT_0</ID>580 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>478</ID>
<type>DE_TO</type>
<position>-8.5,-21</position>
<input>
<ID>IN_0</ID>426 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>801</ID>
<type>DD_KEYPAD_HEX</type>
<position>-81,8.5</position>
<output>
<ID>OUT_0</ID>740 </output>
<output>
<ID>OUT_1</ID>738 </output>
<output>
<ID>OUT_2</ID>739 </output>
<output>
<ID>OUT_3</ID>737 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>479</ID>
<type>DA_FROM</type>
<position>24,-4</position>
<input>
<ID>IN_0</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr1</lparam></gate>
<gate>
<ID>810</ID>
<type>DE_TO</type>
<position>-25,24</position>
<input>
<ID>IN_0</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr8</lparam></gate>
<gate>
<ID>657</ID>
<type>DA_FROM</type>
<position>116,-38</position>
<input>
<ID>IN_0</ID>587 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr10</lparam></gate>
<gate>
<ID>480</ID>
<type>DE_TO</type>
<position>-8.5,-19</position>
<input>
<ID>IN_0</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>481</ID>
<type>DA_FROM</type>
<position>24,4</position>
<input>
<ID>IN_0</ID>459 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>482</ID>
<type>DA_FROM</type>
<position>-38.5,-23.5</position>
<input>
<ID>IN_0</ID>423 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>519</ID>
<type>DA_FROM</type>
<position>43,9.5</position>
<input>
<ID>IN_0</ID>450 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>483</ID>
<type>AI_MUX_8x1</type>
<position>42.5,23</position>
<input>
<ID>IN_0</ID>408 </input>
<input>
<ID>IN_1</ID>439 </input>
<input>
<ID>IN_2</ID>440 </input>
<input>
<ID>IN_3</ID>441 </input>
<input>
<ID>IN_4</ID>431 </input>
<input>
<ID>IN_5</ID>443 </input>
<input>
<ID>IN_6</ID>444 </input>
<input>
<ID>IN_7</ID>445 </input>
<output>
<ID>OUT</ID>446 </output>
<input>
<ID>SEL_0</ID>434 </input>
<input>
<ID>SEL_1</ID>435 </input>
<input>
<ID>SEL_2</ID>436 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>526</ID>
<type>DA_FROM</type>
<position>45,-18.5</position>
<input>
<ID>IN_0</ID>464 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>814</ID>
<type>EE_VDD</type>
<position>-45,23.5</position>
<output>
<ID>OUT_0</ID>745 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>661</ID>
<type>DA_FROM</type>
<position>115.5,24</position>
<input>
<ID>IN_0</ID>562 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>484</ID>
<type>AA_AND2</type>
<position>31,14.5</position>
<input>
<ID>IN_0</ID>438 </input>
<input>
<ID>IN_1</ID>437 </input>
<output>
<ID>OUT</ID>408 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>485</ID>
<type>DA_FROM</type>
<position>24,-10</position>
<input>
<ID>IN_0</ID>452 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr1</lparam></gate>
<gate>
<ID>635</ID>
<type>DE_TO</type>
<position>-14.5,-58</position>
<input>
<ID>IN_0</ID>723 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum3</lparam></gate>
<gate>
<ID>486</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-81,-50</position>
<input>
<ID>IN_0</ID>678 </input>
<input>
<ID>IN_1</ID>679 </input>
<input>
<ID>IN_2</ID>680 </input>
<input>
<ID>IN_3</ID>681 </input>
<input>
<ID>IN_B_0</ID>685 </input>
<input>
<ID>IN_B_1</ID>684 </input>
<input>
<ID>IN_B_2</ID>683 </input>
<input>
<ID>IN_B_3</ID>682 </input>
<output>
<ID>OUT_0</ID>711 </output>
<output>
<ID>OUT_1</ID>712 </output>
<output>
<ID>OUT_2</ID>714 </output>
<output>
<ID>OUT_3</ID>713 </output>
<input>
<ID>carry_in</ID>430 </input>
<output>
<ID>carry_out</ID>621 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>809</ID>
<type>DE_TO</type>
<position>-25,28</position>
<input>
<ID>IN_0</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr10</lparam></gate>
<gate>
<ID>487</ID>
<type>FF_GND</type>
<position>36,-25.5</position>
<output>
<ID>OUT_0</ID>475 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>514</ID>
<type>AA_AND2</type>
<position>31.5,-9.5</position>
<input>
<ID>IN_0</ID>453 </input>
<input>
<ID>IN_1</ID>452 </input>
<output>
<ID>OUT</ID>447 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>665</ID>
<type>DA_FROM</type>
<position>136.5,33.5</position>
<input>
<ID>IN_0</ID>554 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>488</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-34,-50</position>
<input>
<ID>IN_0</ID>697 </input>
<input>
<ID>IN_1</ID>696 </input>
<input>
<ID>IN_2</ID>695 </input>
<input>
<ID>IN_3</ID>694 </input>
<input>
<ID>IN_B_0</ID>701 </input>
<input>
<ID>IN_B_1</ID>700 </input>
<input>
<ID>IN_B_2</ID>699 </input>
<input>
<ID>IN_B_3</ID>698 </input>
<output>
<ID>OUT_0</ID>722 </output>
<output>
<ID>OUT_1</ID>721 </output>
<output>
<ID>OUT_2</ID>720 </output>
<output>
<ID>OUT_3</ID>719 </output>
<input>
<ID>carry_in</ID>428 </input>
<output>
<ID>carry_out</ID>429 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>489</ID>
<type>AI_MUX_8x1</type>
<position>43,-29</position>
<input>
<ID>IN_0</ID>462 </input>
<input>
<ID>IN_1</ID>469 </input>
<input>
<ID>IN_2</ID>470 </input>
<input>
<ID>IN_3</ID>415 </input>
<input>
<ID>IN_4</ID>463 </input>
<input>
<ID>IN_5</ID>473 </input>
<input>
<ID>IN_6</ID>474 </input>
<input>
<ID>IN_7</ID>475 </input>
<output>
<ID>OUT</ID>476 </output>
<input>
<ID>SEL_0</ID>464 </input>
<input>
<ID>SEL_1</ID>465 </input>
<input>
<ID>SEL_2</ID>466 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>490</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-11.5,-50</position>
<input>
<ID>IN_0</ID>705 </input>
<input>
<ID>IN_1</ID>704 </input>
<input>
<ID>IN_2</ID>703 </input>
<input>
<ID>IN_3</ID>702 </input>
<input>
<ID>IN_B_0</ID>709 </input>
<input>
<ID>IN_B_1</ID>708 </input>
<input>
<ID>IN_B_2</ID>707 </input>
<input>
<ID>IN_B_3</ID>706 </input>
<output>
<ID>OUT_0</ID>726 </output>
<output>
<ID>OUT_1</ID>725 </output>
<output>
<ID>OUT_2</ID>724 </output>
<output>
<ID>OUT_3</ID>723 </output>
<input>
<ID>carry_in</ID>710 </input>
<output>
<ID>carry_out</ID>428 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>527</ID>
<type>DA_FROM</type>
<position>41,-18.5</position>
<input>
<ID>IN_0</ID>466 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>491</ID>
<type>AE_SMALL_INVERTER</type>
<position>31.5,-28</position>
<input>
<ID>IN_0</ID>472 </input>
<output>
<ID>OUT_0</ID>463 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>669</ID>
<type>AA_AND2</type>
<position>123.5,-9.5</position>
<input>
<ID>IN_0</ID>573 </input>
<input>
<ID>IN_1</ID>572 </input>
<output>
<ID>OUT</ID>567 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>492</ID>
<type>AE_SMALL_INVERTER</type>
<position>31,24</position>
<input>
<ID>IN_0</ID>442 </input>
<output>
<ID>OUT_0</ID>431 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>493</ID>
<type>DA_FROM</type>
<position>24,-32</position>
<input>
<ID>IN_0</ID>470 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr2</lparam></gate>
<gate>
<ID>494</ID>
<type>DA_FROM</type>
<position>23.5,18</position>
<input>
<ID>IN_0</ID>439 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum0</lparam></gate>
<gate>
<ID>515</ID>
<type>DA_FROM</type>
<position>24,2</position>
<input>
<ID>IN_0</ID>458 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>522</ID>
<type>AA_AND2</type>
<position>31.5,-37.5</position>
<input>
<ID>IN_0</ID>468 </input>
<input>
<ID>IN_1</ID>467 </input>
<output>
<ID>OUT</ID>462 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>495</ID>
<type>DA_FROM</type>
<position>24,-26</position>
<input>
<ID>IN_0</ID>473 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>817</ID>
<type>BW_8X1_BUS_END</type>
<position>-31.5,12</position>
<input>
<ID>IN_0</ID>734 </input>
<input>
<ID>IN_1</ID>733 </input>
<input>
<ID>IN_2</ID>732 </input>
<input>
<ID>IN_3</ID>731 </input>
<input>
<ID>IN_4</ID>730 </input>
<input>
<ID>IN_5</ID>729 </input>
<input>
<ID>IN_6</ID>728 </input>
<input>
<ID>IN_7</ID>727 </input>
<input>
<ID>OUT</ID>651 652 653 654 655 656 657 658 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>496</ID>
<type>DA_FROM</type>
<position>23.5,20</position>
<input>
<ID>IN_0</ID>440 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr0</lparam></gate>
<gate>
<ID>673</ID>
<type>DA_FROM</type>
<position>116,-8</position>
<input>
<ID>IN_0</ID>573 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>512</ID>
<type>DA_FROM</type>
<position>42.5,33.5</position>
<input>
<ID>IN_0</ID>435 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>497</ID>
<type>DA_FROM</type>
<position>24,-28</position>
<input>
<ID>IN_0</ID>472 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>704</ID>
<type>DA_FROM</type>
<position>159,19.5</position>
<input>
<ID>IN_0</ID>620 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr12</lparam></gate>
<gate>
<ID>498</ID>
<type>DA_FROM</type>
<position>23.5,28</position>
<input>
<ID>IN_0</ID>444 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>535</ID>
<type>DA_FROM</type>
<position>25,-53</position>
<input>
<ID>IN_0</ID>488 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>499</ID>
<type>DA_FROM</type>
<position>24,-38</position>
<input>
<ID>IN_0</ID>467 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr2</lparam></gate>
<gate>
<ID>500</ID>
<type>DA_FROM</type>
<position>23.5,26</position>
<input>
<ID>IN_0</ID>443 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>677</ID>
<type>DA_FROM</type>
<position>133,9.5</position>
<input>
<ID>IN_0</ID>571 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>516</ID>
<type>DA_FROM</type>
<position>24,0</position>
<input>
<ID>IN_0</ID>457 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>501</ID>
<type>DA_FROM</type>
<position>43,-18.5</position>
<input>
<ID>IN_0</ID>465 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>708</ID>
<type>DA_FROM</type>
<position>117,-65</position>
<input>
<ID>IN_0</ID>602 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr11</lparam></gate>
<gate>
<ID>523</ID>
<type>DA_FROM</type>
<position>24,-34</position>
<input>
<ID>IN_0</ID>469 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum2</lparam></gate>
<gate>
<ID>502</ID>
<type>DA_FROM</type>
<position>23.5,22</position>
<input>
<ID>IN_0</ID>441 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr0</lparam></gate>
<gate>
<ID>503</ID>
<type>FF_GND</type>
<position>37,-52.5</position>
<output>
<ID>OUT_0</ID>490 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>504</ID>
<type>CC_PRI_ENCODER_8x3</type>
<position>-20,-17</position>
<input>
<ID>ENABLE</ID>424 </input>
<input>
<ID>IN_0</ID>423 </input>
<input>
<ID>IN_1</ID>422 </input>
<input>
<ID>IN_2</ID>421 </input>
<input>
<ID>IN_3</ID>420 </input>
<input>
<ID>IN_4</ID>419 </input>
<input>
<ID>IN_5</ID>418 </input>
<input>
<ID>IN_6</ID>417 </input>
<input>
<ID>IN_7</ID>416 </input>
<output>
<ID>OUT_0</ID>427 </output>
<output>
<ID>OUT_1</ID>426 </output>
<output>
<ID>OUT_2</ID>425 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>681</ID>
<type>DE_TO</type>
<position>183.5,-1.5</position>
<input>
<ID>IN_0</ID>641 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin13</lparam></gate>
<gate>
<ID>520</ID>
<type>DA_FROM</type>
<position>41,9.5</position>
<input>
<ID>IN_0</ID>451 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>505</ID>
<type>FF_GND</type>
<position>-38,-9.5</position>
<output>
<ID>OUT_0</ID>416 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>712</ID>
<type>AI_MUX_8x1</type>
<position>178.5,-1.5</position>
<input>
<ID>IN_0</ID>627 </input>
<input>
<ID>IN_1</ID>634 </input>
<input>
<ID>IN_2</ID>635 </input>
<input>
<ID>IN_3</ID>576 </input>
<input>
<ID>IN_4</ID>628 </input>
<input>
<ID>IN_5</ID>638 </input>
<input>
<ID>IN_6</ID>639 </input>
<input>
<ID>IN_7</ID>640 </input>
<output>
<ID>OUT</ID>641 </output>
<input>
<ID>SEL_0</ID>629 </input>
<input>
<ID>SEL_1</ID>630 </input>
<input>
<ID>SEL_2</ID>631 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>506</ID>
<type>EE_VDD</type>
<position>-24,-9.5</position>
<output>
<ID>OUT_0</ID>424 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>543</ID>
<type>DA_FROM</type>
<position>159.5,1.5</position>
<input>
<ID>IN_0</ID>638 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>507</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-57.5,-50</position>
<input>
<ID>IN_0</ID>688 </input>
<input>
<ID>IN_1</ID>689 </input>
<input>
<ID>IN_2</ID>687 </input>
<input>
<ID>IN_3</ID>686 </input>
<input>
<ID>IN_B_0</ID>693 </input>
<input>
<ID>IN_B_1</ID>692 </input>
<input>
<ID>IN_B_2</ID>691 </input>
<input>
<ID>IN_B_3</ID>690 </input>
<output>
<ID>OUT_0</ID>718 </output>
<output>
<ID>OUT_1</ID>717 </output>
<output>
<ID>OUT_2</ID>716 </output>
<output>
<ID>OUT_3</ID>715 </output>
<input>
<ID>carry_in</ID>429 </input>
<output>
<ID>carry_out</ID>430 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>508</ID>
<type>DA_FROM</type>
<position>23.5,24</position>
<input>
<ID>IN_0</ID>442 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>685</ID>
<type>BV_4x1_BUS_END</type>
<position>-50,10</position>
<input>
<ID>IN_0</ID>399 </input>
<input>
<ID>IN_1</ID>401 </input>
<input>
<ID>IN_2</ID>398 </input>
<input>
<ID>IN_3</ID>400 </input>
<input>
<ID>OUT</ID>750 751 752 753 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>524</ID>
<type>DA_FROM</type>
<position>24,-24</position>
<input>
<ID>IN_0</ID>474 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>509</ID>
<type>DA_FROM</type>
<position>23.5,16</position>
<input>
<ID>IN_0</ID>438 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>716</ID>
<type>FF_GND</type>
<position>171.5,-26</position>
<output>
<ID>OUT_0</ID>662 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>510</ID>
<type>DA_FROM</type>
<position>23.5,14</position>
<input>
<ID>IN_0</ID>437 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr0</lparam></gate>
<gate>
<ID>531</ID>
<type>AE_SMALL_INVERTER</type>
<position>32.5,-55</position>
<input>
<ID>IN_0</ID>487 </input>
<output>
<ID>OUT_0</ID>478 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>511</ID>
<type>DA_FROM</type>
<position>44.5,33.5</position>
<input>
<ID>IN_0</ID>434 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>528</ID>
<type>DE_TO</type>
<position>49,-56</position>
<input>
<ID>IN_0</ID>491 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin3</lparam></gate>
<gate>
<ID>529</ID>
<type>AI_MUX_8x1</type>
<position>44,-56</position>
<input>
<ID>IN_0</ID>477 </input>
<input>
<ID>IN_1</ID>484 </input>
<input>
<ID>IN_2</ID>485 </input>
<input>
<ID>IN_3</ID>432 </input>
<input>
<ID>IN_4</ID>478 </input>
<input>
<ID>IN_5</ID>488 </input>
<input>
<ID>IN_6</ID>489 </input>
<input>
<ID>IN_7</ID>490 </input>
<output>
<ID>OUT</ID>491 </output>
<input>
<ID>SEL_0</ID>479 </input>
<input>
<ID>SEL_1</ID>480 </input>
<input>
<ID>SEL_2</ID>481 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>530</ID>
<type>AA_AND2</type>
<position>32.5,-64.5</position>
<input>
<ID>IN_0</ID>483 </input>
<input>
<ID>IN_1</ID>482 </input>
<output>
<ID>OUT</ID>477 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>532</ID>
<type>DA_FROM</type>
<position>25,-61</position>
<input>
<ID>IN_0</ID>484 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum3</lparam></gate>
<gate>
<ID>533</ID>
<type>DA_FROM</type>
<position>25,-59</position>
<input>
<ID>IN_0</ID>485 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr3</lparam></gate>
<gate>
<ID>534</ID>
<type>DA_FROM</type>
<position>25,-51</position>
<input>
<ID>IN_0</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>536</ID>
<type>DA_FROM</type>
<position>25,-55</position>
<input>
<ID>IN_0</ID>487 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>537</ID>
<type>DA_FROM</type>
<position>25,-63</position>
<input>
<ID>IN_0</ID>483 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>538</ID>
<type>DA_FROM</type>
<position>25,-65</position>
<input>
<ID>IN_0</ID>482 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr3</lparam></gate>
<gate>
<ID>539</ID>
<type>DA_FROM</type>
<position>46,-45.5</position>
<input>
<ID>IN_0</ID>479 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>540</ID>
<type>DA_FROM</type>
<position>159,25.5</position>
<input>
<ID>IN_0</ID>623 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>541</ID>
<type>DA_FROM</type>
<position>44,-45.5</position>
<input>
<ID>IN_0</ID>480 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>542</ID>
<type>DA_FROM</type>
<position>42,-45.5</position>
<input>
<ID>IN_0</ID>481 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>544</ID>
<type>FF_GND</type>
<position>83,26.5</position>
<output>
<ID>OUT_0</ID>505 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>545</ID>
<type>DE_TO</type>
<position>95,23</position>
<input>
<ID>IN_0</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin4</lparam></gate>
<gate>
<ID>546</ID>
<type>DA_FROM</type>
<position>159,15.5</position>
<input>
<ID>IN_0</ID>618 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>547</ID>
<type>FF_GND</type>
<position>83.5,2.5</position>
<output>
<ID>OUT_0</ID>520 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>548</ID>
<type>DE_TO</type>
<position>95.5,-1</position>
<input>
<ID>IN_0</ID>521 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin5</lparam></gate>
<gate>
<ID>549</ID>
<type>DA_FROM</type>
<position>159,27.5</position>
<input>
<ID>IN_0</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>550</ID>
<type>AI_MUX_8x1</type>
<position>90.5,-1</position>
<input>
<ID>IN_0</ID>507 </input>
<input>
<ID>IN_1</ID>514 </input>
<input>
<ID>IN_2</ID>515 </input>
<input>
<ID>IN_3</ID>456 </input>
<input>
<ID>IN_4</ID>508 </input>
<input>
<ID>IN_5</ID>518 </input>
<input>
<ID>IN_6</ID>519 </input>
<input>
<ID>IN_7</ID>520 </input>
<output>
<ID>OUT</ID>521 </output>
<input>
<ID>SEL_0</ID>509 </input>
<input>
<ID>SEL_1</ID>510 </input>
<input>
<ID>SEL_2</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>551</ID>
<type>AE_SMALL_INVERTER</type>
<position>79,0</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>508 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>552</ID>
<type>DA_FROM</type>
<position>176,33</position>
<input>
<ID>IN_0</ID>616 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>553</ID>
<type>DA_FROM</type>
<position>71.5,-6</position>
<input>
<ID>IN_0</ID>514 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum5</lparam></gate>
<gate>
<ID>554</ID>
<type>DA_FROM</type>
<position>71.5,-4</position>
<input>
<ID>IN_0</ID>515 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr5</lparam></gate>
<gate>
<ID>555</ID>
<type>AA_AND2</type>
<position>167,-38</position>
<input>
<ID>IN_0</ID>648 </input>
<input>
<ID>IN_1</ID>647 </input>
<output>
<ID>OUT</ID>642 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>556</ID>
<type>DA_FROM</type>
<position>71.5,4</position>
<input>
<ID>IN_0</ID>519 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>557</ID>
<type>AI_MUX_8x1</type>
<position>90,23</position>
<input>
<ID>IN_0</ID>492 </input>
<input>
<ID>IN_1</ID>499 </input>
<input>
<ID>IN_2</ID>500 </input>
<input>
<ID>IN_3</ID>433 </input>
<input>
<ID>IN_4</ID>493 </input>
<input>
<ID>IN_5</ID>503 </input>
<input>
<ID>IN_6</ID>504 </input>
<input>
<ID>IN_7</ID>505 </input>
<output>
<ID>OUT</ID>506 </output>
<input>
<ID>SEL_0</ID>494 </input>
<input>
<ID>SEL_1</ID>495 </input>
<input>
<ID>SEL_2</ID>496 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>558</ID>
<type>DA_FROM</type>
<position>159.5,-0.5</position>
<input>
<ID>IN_0</ID>637 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>559</ID>
<type>AA_AND2</type>
<position>78.5,14.5</position>
<input>
<ID>IN_0</ID>498 </input>
<input>
<ID>IN_1</ID>497 </input>
<output>
<ID>OUT</ID>492 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>560</ID>
<type>DA_FROM</type>
<position>71.5,-10</position>
<input>
<ID>IN_0</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr5</lparam></gate>
<gate>
<ID>561</ID>
<type>DA_FROM</type>
<position>180,33</position>
<input>
<ID>IN_0</ID>614 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>562</ID>
<type>FF_GND</type>
<position>83.5,-25.5</position>
<output>
<ID>OUT_0</ID>535 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>563</ID>
<type>AI_MUX_8x1</type>
<position>90.5,-29</position>
<input>
<ID>IN_0</ID>522 </input>
<input>
<ID>IN_1</ID>529 </input>
<input>
<ID>IN_2</ID>530 </input>
<input>
<ID>IN_3</ID>471 </input>
<input>
<ID>IN_4</ID>523 </input>
<input>
<ID>IN_5</ID>533 </input>
<input>
<ID>IN_6</ID>534 </input>
<input>
<ID>IN_7</ID>535 </input>
<output>
<ID>OUT</ID>536 </output>
<input>
<ID>SEL_0</ID>524 </input>
<input>
<ID>SEL_1</ID>525 </input>
<input>
<ID>SEL_2</ID>526 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>564</ID>
<type>DA_FROM</type>
<position>176.5,9</position>
<input>
<ID>IN_0</ID>631 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>565</ID>
<type>AE_SMALL_INVERTER</type>
<position>79,-28</position>
<input>
<ID>IN_0</ID>532 </input>
<output>
<ID>OUT_0</ID>523 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>566</ID>
<type>AE_SMALL_INVERTER</type>
<position>78.5,24</position>
<input>
<ID>IN_0</ID>502 </input>
<output>
<ID>OUT_0</ID>493 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>567</ID>
<type>DE_TO</type>
<position>184.5,-56.5</position>
<input>
<ID>IN_0</ID>677 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin15</lparam></gate>
<gate>
<ID>568</ID>
<type>DA_FROM</type>
<position>71.5,-32</position>
<input>
<ID>IN_0</ID>530 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr6</lparam></gate>
<gate>
<ID>569</ID>
<type>DA_FROM</type>
<position>71,18</position>
<input>
<ID>IN_0</ID>499 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum4</lparam></gate>
<gate>
<ID>570</ID>
<type>DA_FROM</type>
<position>159.5,-24.5</position>
<input>
<ID>IN_0</ID>661 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>571</ID>
<type>DA_FROM</type>
<position>71.5,-26</position>
<input>
<ID>IN_0</ID>533 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>572</ID>
<type>DA_FROM</type>
<position>71,20</position>
<input>
<ID>IN_0</ID>500 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr4</lparam></gate>
<gate>
<ID>573</ID>
<type>DA_FROM</type>
<position>180.5,9</position>
<input>
<ID>IN_0</ID>629 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>574</ID>
<type>DA_FROM</type>
<position>71.5,-28</position>
<input>
<ID>IN_0</ID>532 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>575</ID>
<type>DA_FROM</type>
<position>71,28</position>
<input>
<ID>IN_0</ID>504 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>576</ID>
<type>DA_FROM</type>
<position>176.5,-19</position>
<input>
<ID>IN_0</ID>646 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>577</ID>
<type>DA_FROM</type>
<position>71.5,-38</position>
<input>
<ID>IN_0</ID>527 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr6</lparam></gate>
<gate>
<ID>578</ID>
<type>DA_FROM</type>
<position>71,26</position>
<input>
<ID>IN_0</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>579</ID>
<type>DA_FROM</type>
<position>90.5,-18.5</position>
<input>
<ID>IN_0</ID>525 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>580</ID>
<type>DE_TO</type>
<position>-25,32</position>
<input>
<ID>IN_0</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr12</lparam></gate>
<gate>
<ID>581</ID>
<type>AA_AND2</type>
<position>168,-65</position>
<input>
<ID>IN_0</ID>670 </input>
<input>
<ID>IN_1</ID>669 </input>
<output>
<ID>OUT</ID>664 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>582</ID>
<type>DA_FROM</type>
<position>71,24</position>
<input>
<ID>IN_0</ID>502 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>583</ID>
<type>DA_FROM</type>
<position>71,16</position>
<input>
<ID>IN_0</ID>498 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>584</ID>
<type>DA_FROM</type>
<position>159.5,-36.5</position>
<input>
<ID>IN_0</ID>648 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>585</ID>
<type>DA_FROM</type>
<position>71,14</position>
<input>
<ID>IN_0</ID>497 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr4</lparam></gate>
<gate>
<ID>586</ID>
<type>DA_FROM</type>
<position>92,33.5</position>
<input>
<ID>IN_0</ID>494 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>587</ID>
<type>DA_FROM</type>
<position>160.5,-51.5</position>
<input>
<ID>IN_0</ID>675 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>588</ID>
<type>DA_FROM</type>
<position>90,33.5</position>
<input>
<ID>IN_0</ID>495 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>589</ID>
<type>DA_FROM</type>
<position>88,33.5</position>
<input>
<ID>IN_0</ID>496 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>590</ID>
<type>AA_AND2</type>
<position>79,-9.5</position>
<input>
<ID>IN_0</ID>513 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>507 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>591</ID>
<type>DA_FROM</type>
<position>71.5,2</position>
<input>
<ID>IN_0</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>592</ID>
<type>DA_FROM</type>
<position>160.5,-63.5</position>
<input>
<ID>IN_0</ID>670 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>593</ID>
<type>BV_4x1_BUS_END</type>
<position>-71.5,-6</position>
<input>
<ID>IN_0</ID>744 </input>
<input>
<ID>IN_1</ID>743 </input>
<input>
<ID>IN_2</ID>742 </input>
<input>
<ID>IN_3</ID>741 </input>
<input>
<ID>OUT</ID>750 751 752 753 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>594</ID>
<type>DA_FROM</type>
<position>71.5,0</position>
<input>
<ID>IN_0</ID>517 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>595</ID>
<type>DA_FROM</type>
<position>160.5,-61.5</position>
<input>
<ID>IN_0</ID>671 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum15</lparam></gate>
<gate>
<ID>596</ID>
<type>DA_FROM</type>
<position>71.5,-8</position>
<input>
<ID>IN_0</ID>513 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>597</ID>
<type>DA_FROM</type>
<position>92.5,9.5</position>
<input>
<ID>IN_0</ID>509 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>598</ID>
<type>DA_FROM</type>
<position>90.5,9.5</position>
<input>
<ID>IN_0</ID>510 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>599</ID>
<type>DA_FROM</type>
<position>88.5,9.5</position>
<input>
<ID>IN_0</ID>511 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>600</ID>
<type>DE_TO</type>
<position>95.5,-29</position>
<input>
<ID>IN_0</ID>536 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin6</lparam></gate>
<gate>
<ID>601</ID>
<type>AA_AND2</type>
<position>79,-37.5</position>
<input>
<ID>IN_0</ID>528 </input>
<input>
<ID>IN_1</ID>527 </input>
<output>
<ID>OUT</ID>522 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>602</ID>
<type>DA_FROM</type>
<position>71.5,-34</position>
<input>
<ID>IN_0</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum6</lparam></gate>
<gate>
<ID>603</ID>
<type>DA_FROM</type>
<position>71.5,-24</position>
<input>
<ID>IN_0</ID>534 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>604</ID>
<type>DA_FROM</type>
<position>71.5,-36</position>
<input>
<ID>IN_0</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>605</ID>
<type>DA_FROM</type>
<position>92.5,-18.5</position>
<input>
<ID>IN_0</ID>524 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>606</ID>
<type>DA_FROM</type>
<position>88.5,-18.5</position>
<input>
<ID>IN_0</ID>526 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>607</ID>
<type>FF_GND</type>
<position>84.5,-52.5</position>
<output>
<ID>OUT_0</ID>550 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>608</ID>
<type>DE_TO</type>
<position>96.5,-56</position>
<input>
<ID>IN_0</ID>551 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin7</lparam></gate>
<gate>
<ID>609</ID>
<type>AI_MUX_8x1</type>
<position>91.5,-56</position>
<input>
<ID>IN_0</ID>537 </input>
<input>
<ID>IN_1</ID>544 </input>
<input>
<ID>IN_2</ID>545 </input>
<input>
<ID>IN_3</ID>486 </input>
<input>
<ID>IN_4</ID>538 </input>
<input>
<ID>IN_5</ID>548 </input>
<input>
<ID>IN_6</ID>549 </input>
<input>
<ID>IN_7</ID>550 </input>
<output>
<ID>OUT</ID>551 </output>
<input>
<ID>SEL_0</ID>539 </input>
<input>
<ID>SEL_1</ID>540 </input>
<input>
<ID>SEL_2</ID>541 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>610</ID>
<type>AA_AND2</type>
<position>80,-64.5</position>
<input>
<ID>IN_0</ID>543 </input>
<input>
<ID>IN_1</ID>542 </input>
<output>
<ID>OUT</ID>537 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>611</ID>
<type>AE_SMALL_INVERTER</type>
<position>80,-55</position>
<input>
<ID>IN_0</ID>547 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>612</ID>
<type>DA_FROM</type>
<position>72.5,-61</position>
<input>
<ID>IN_0</ID>544 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum7</lparam></gate>
<gate>
<ID>613</ID>
<type>DA_FROM</type>
<position>72.5,-59</position>
<input>
<ID>IN_0</ID>545 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr7</lparam></gate>
<gate>
<ID>614</ID>
<type>DA_FROM</type>
<position>72.5,-51</position>
<input>
<ID>IN_0</ID>549 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>615</ID>
<type>DA_FROM</type>
<position>72.5,-53</position>
<input>
<ID>IN_0</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>616</ID>
<type>DA_FROM</type>
<position>72.5,-55</position>
<input>
<ID>IN_0</ID>547 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>617</ID>
<type>DA_FROM</type>
<position>72.5,-63</position>
<input>
<ID>IN_0</ID>543 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>618</ID>
<type>DA_FROM</type>
<position>72.5,-65</position>
<input>
<ID>IN_0</ID>542 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr7</lparam></gate>
<gate>
<ID>620</ID>
<type>DA_FROM</type>
<position>-36.5,-38</position>
<input>
<ID>IN_0</ID>696 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>621</ID>
<type>DA_FROM</type>
<position>91.5,-45.5</position>
<input>
<ID>IN_0</ID>540 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>622</ID>
<type>DA_FROM</type>
<position>89.5,-45.5</position>
<input>
<ID>IN_0</ID>541 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>623</ID>
<type>DA_FROM</type>
<position>-87.5,-38.5</position>
<input>
<ID>IN_0</ID>681 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>991</ID>
<type>AA_LABEL</type>
<position>-69,53.5</position>
<gparam>LABEL_TEXT ALU</gparam>
<gparam>TEXT_HEIGHT 10</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>624</ID>
<type>FF_GND</type>
<position>127.5,26.5</position>
<output>
<ID>OUT_0</ID>565 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>625</ID>
<type>DE_TO</type>
<position>139.5,23</position>
<input>
<ID>IN_0</ID>566 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin8</lparam></gate>
<gate>
<ID>626</ID>
<type>DA_FROM</type>
<position>-61,-38</position>
<input>
<ID>IN_0</ID>689 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>628</ID>
<type>DE_TO</type>
<position>140,-1</position>
<input>
<ID>IN_0</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin9</lparam></gate>
<gate>
<ID>629</ID>
<type>DA_FROM</type>
<position>-19,-38</position>
<input>
<ID>IN_0</ID>702 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>630</ID>
<type>AI_MUX_8x1</type>
<position>135,-1</position>
<input>
<ID>IN_0</ID>567 </input>
<input>
<ID>IN_1</ID>574 </input>
<input>
<ID>IN_2</ID>575 </input>
<input>
<ID>IN_3</ID>516 </input>
<input>
<ID>IN_4</ID>568 </input>
<input>
<ID>IN_5</ID>578 </input>
<input>
<ID>IN_6</ID>579 </input>
<input>
<ID>IN_7</ID>580 </input>
<output>
<ID>OUT</ID>581 </output>
<input>
<ID>SEL_0</ID>569 </input>
<input>
<ID>SEL_1</ID>570 </input>
<input>
<ID>SEL_2</ID>571 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>632</ID>
<type>DA_FROM</type>
<position>-83.5,-38.5</position>
<input>
<ID>IN_0</ID>679 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>633</ID>
<type>DA_FROM</type>
<position>116,-6</position>
<input>
<ID>IN_0</ID>574 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum9</lparam></gate>
<gate>
<ID>634</ID>
<type>DA_FROM</type>
<position>116,-4</position>
<input>
<ID>IN_0</ID>575 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr9</lparam></gate>
<gate>
<ID>636</ID>
<type>DA_FROM</type>
<position>116,4</position>
<input>
<ID>IN_0</ID>579 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>637</ID>
<type>AI_MUX_8x1</type>
<position>134.5,23</position>
<input>
<ID>IN_0</ID>552 </input>
<input>
<ID>IN_1</ID>559 </input>
<input>
<ID>IN_2</ID>560 </input>
<input>
<ID>IN_3</ID>501 </input>
<input>
<ID>IN_4</ID>553 </input>
<input>
<ID>IN_5</ID>563 </input>
<input>
<ID>IN_6</ID>564 </input>
<input>
<ID>IN_7</ID>565 </input>
<output>
<ID>OUT</ID>566 </output>
<input>
<ID>SEL_0</ID>554 </input>
<input>
<ID>SEL_1</ID>555 </input>
<input>
<ID>SEL_2</ID>556 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>638</ID>
<type>FF_GND</type>
<position>-2,-50.5</position>
<output>
<ID>OUT_0</ID>710 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>640</ID>
<type>DA_FROM</type>
<position>116,-10</position>
<input>
<ID>IN_0</ID>572 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr9</lparam></gate>
<gate>
<ID>642</ID>
<type>FF_GND</type>
<position>128,-25.5</position>
<output>
<ID>OUT_0</ID>595 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>643</ID>
<type>AI_MUX_8x1</type>
<position>135,-29</position>
<input>
<ID>IN_0</ID>582 </input>
<input>
<ID>IN_1</ID>589 </input>
<input>
<ID>IN_2</ID>590 </input>
<input>
<ID>IN_3</ID>531 </input>
<input>
<ID>IN_4</ID>583 </input>
<input>
<ID>IN_5</ID>593 </input>
<input>
<ID>IN_6</ID>594 </input>
<input>
<ID>IN_7</ID>595 </input>
<output>
<ID>OUT</ID>596 </output>
<input>
<ID>SEL_0</ID>584 </input>
<input>
<ID>SEL_1</ID>585 </input>
<input>
<ID>SEL_2</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>804</ID>
<type>AE_REGISTER8</type>
<position>-44,11.5</position>
<input>
<ID>IN_0</ID>399 </input>
<input>
<ID>IN_1</ID>401 </input>
<input>
<ID>IN_2</ID>398 </input>
<input>
<ID>IN_3</ID>400 </input>
<input>
<ID>IN_4</ID>402 </input>
<input>
<ID>IN_5</ID>403 </input>
<input>
<ID>IN_6</ID>404 </input>
<input>
<ID>IN_7</ID>405 </input>
<output>
<ID>OUT_0</ID>636 </output>
<output>
<ID>OUT_1</ID>411 </output>
<output>
<ID>OUT_2</ID>406 </output>
<output>
<ID>OUT_3</ID>412 </output>
<output>
<ID>OUT_4</ID>409 </output>
<output>
<ID>OUT_5</ID>413 </output>
<output>
<ID>OUT_6</ID>407 </output>
<output>
<ID>OUT_7</ID>410 </output>
<input>
<ID>clock</ID>735 </input>
<input>
<ID>count_enable</ID>736 </input>
<input>
<ID>load</ID>745 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 106</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>644</ID>
<type>DE_TO</type>
<position>-10.5,-58</position>
<input>
<ID>IN_0</ID>725 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum1</lparam></gate>
<gate>
<ID>646</ID>
<type>AE_SMALL_INVERTER</type>
<position>123,24</position>
<input>
<ID>IN_0</ID>562 </input>
<output>
<ID>OUT_0</ID>553 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>647</ID>
<type>DE_TO</type>
<position>-60.5,-58.5</position>
<input>
<ID>IN_0</ID>715 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum11</lparam></gate>
<gate>
<ID>792</ID>
<type>DA_FROM</type>
<position>116,-2</position>
<input>
<ID>IN_0</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr9</lparam></gate>
<gate>
<ID>648</ID>
<type>DA_FROM</type>
<position>116,-32</position>
<input>
<ID>IN_0</ID>590 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr10</lparam></gate>
<gate>
<ID>650</ID>
<type>DE_TO</type>
<position>-33,-58.5</position>
<input>
<ID>IN_0</ID>721 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum5</lparam></gate>
<gate>
<ID>651</ID>
<type>DA_FROM</type>
<position>116,-26</position>
<input>
<ID>IN_0</ID>593 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>812</ID>
<type>BV_4x1_BUS_END</type>
<position>-50,22</position>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>652</ID>
<type>DA_FROM</type>
<position>115.5,20</position>
<input>
<ID>IN_0</ID>560 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr8</lparam></gate>
<gate>
<ID>654</ID>
<type>DA_FROM</type>
<position>116,-28</position>
<input>
<ID>IN_0</ID>592 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>655</ID>
<type>DA_FROM</type>
<position>115.5,28</position>
<input>
<ID>IN_0</ID>564 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>800</ID>
<type>DD_KEYPAD_HEX</type>
<position>-81,-6</position>
<output>
<ID>OUT_0</ID>744 </output>
<output>
<ID>OUT_1</ID>743 </output>
<output>
<ID>OUT_2</ID>742 </output>
<output>
<ID>OUT_3</ID>741 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 10</lparam></gate>
<gate>
<ID>656</ID>
<type>DE_TO</type>
<position>-56.5,-58.5</position>
<input>
<ID>IN_0</ID>717 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum9</lparam></gate>
<gate>
<ID>658</ID>
<type>DA_FROM</type>
<position>115.5,26</position>
<input>
<ID>IN_0</ID>563 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>659</ID>
<type>DA_FROM</type>
<position>135,-18.5</position>
<input>
<ID>IN_0</ID>585 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>660</ID>
<type>DE_TO</type>
<position>-80,-58.5</position>
<input>
<ID>IN_0</ID>712 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum13</lparam></gate>
<gate>
<ID>662</ID>
<type>DA_FROM</type>
<position>115.5,16</position>
<input>
<ID>IN_0</ID>558 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>663</ID>
<type>DE_TO</type>
<position>-37,-58.5</position>
<input>
<ID>IN_0</ID>719 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum7</lparam></gate>
<gate>
<ID>808</ID>
<type>DE_TO</type>
<position>-25,30</position>
<input>
<ID>IN_0</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr11</lparam></gate>
<gate>
<ID>664</ID>
<type>DA_FROM</type>
<position>115.5,14</position>
<input>
<ID>IN_0</ID>557 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr8</lparam></gate>
<gate>
<ID>666</ID>
<type>DA_FROM</type>
<position>134.5,33.5</position>
<input>
<ID>IN_0</ID>555 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>667</ID>
<type>DA_FROM</type>
<position>132.5,33.5</position>
<input>
<ID>IN_0</ID>556 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>668</ID>
<type>DE_TO</type>
<position>183,22.5</position>
<input>
<ID>IN_0</ID>626 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin12</lparam></gate>
<gate>
<ID>670</ID>
<type>DA_FROM</type>
<position>116,2</position>
<input>
<ID>IN_0</ID>578 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>671</ID>
<type>DA_FROM</type>
<position>116,0</position>
<input>
<ID>IN_0</ID>577 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>816</ID>
<type>BW_8X1_BUS_END</type>
<position>-38,12</position>
<input>
<ID>IN_0</ID>636 </input>
<input>
<ID>IN_1</ID>411 </input>
<input>
<ID>IN_2</ID>406 </input>
<input>
<ID>IN_3</ID>412 </input>
<input>
<ID>IN_4</ID>409 </input>
<input>
<ID>IN_5</ID>413 </input>
<input>
<ID>IN_6</ID>407 </input>
<input>
<ID>IN_7</ID>410 </input>
<input>
<ID>OUT</ID>651 652 653 654 655 656 657 658 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>672</ID>
<type>DE_TO</type>
<position>-84,-58.5</position>
<input>
<ID>IN_0</ID>713 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum15</lparam></gate>
<gate>
<ID>674</ID>
<type>DA_FROM</type>
<position>137,9.5</position>
<input>
<ID>IN_0</ID>569 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>675</ID>
<type>DA_FROM</type>
<position>134,-45.5</position>
<input>
<ID>IN_0</ID>601 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>676</ID>
<type>DA_FROM</type>
<position>135,9.5</position>
<input>
<ID>IN_0</ID>570 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>678</ID>
<type>AI_MUX_8x1</type>
<position>178,22.5</position>
<input>
<ID>IN_0</ID>612 </input>
<input>
<ID>IN_1</ID>619 </input>
<input>
<ID>IN_2</ID>620 </input>
<input>
<ID>IN_3</ID>561 </input>
<input>
<ID>IN_4</ID>613 </input>
<input>
<ID>IN_5</ID>623 </input>
<input>
<ID>IN_6</ID>624 </input>
<input>
<ID>IN_7</ID>625 </input>
<output>
<ID>OUT</ID>626 </output>
<input>
<ID>SEL_0</ID>614 </input>
<input>
<ID>SEL_1</ID>615 </input>
<input>
<ID>SEL_2</ID>616 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>679</ID>
<type>DE_TO</type>
<position>140,-29</position>
<input>
<ID>IN_0</ID>596 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin10</lparam></gate>
<gate>
<ID>680</ID>
<type>AA_AND2</type>
<position>123.5,-37.5</position>
<input>
<ID>IN_0</ID>588 </input>
<input>
<ID>IN_1</ID>587 </input>
<output>
<ID>OUT</ID>582 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>682</ID>
<type>DA_FROM</type>
<position>116,-34</position>
<input>
<ID>IN_0</ID>589 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum10</lparam></gate>
<gate>
<ID>683</ID>
<type>DA_FROM</type>
<position>116,-24</position>
<input>
<ID>IN_0</ID>594 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>684</ID>
<type>DA_FROM</type>
<position>138,-45.5</position>
<input>
<ID>IN_0</ID>599 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>686</ID>
<type>DA_FROM</type>
<position>116,-36</position>
<input>
<ID>IN_0</ID>588 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>687</ID>
<type>DA_FROM</type>
<position>159.5,-4.5</position>
<input>
<ID>IN_0</ID>635 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr13</lparam></gate>
<gate>
<ID>688</ID>
<type>DA_FROM</type>
<position>137,-18.5</position>
<input>
<ID>IN_0</ID>584 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>689</ID>
<type>DA_FROM</type>
<position>133,-18.5</position>
<input>
<ID>IN_0</ID>586 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>690</ID>
<type>DA_FROM</type>
<position>159,17.5</position>
<input>
<ID>IN_0</ID>619 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum12</lparam></gate>
<gate>
<ID>691</ID>
<type>FF_GND</type>
<position>129,-52.5</position>
<output>
<ID>OUT_0</ID>610 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>692</ID>
<type>DE_TO</type>
<position>141,-56</position>
<input>
<ID>IN_0</ID>611 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin11</lparam></gate>
<gate>
<ID>693</ID>
<type>DA_FROM</type>
<position>159.5,-10.5</position>
<input>
<ID>IN_0</ID>632 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr13</lparam></gate>
<gate>
<ID>694</ID>
<type>AI_MUX_8x1</type>
<position>136,-56</position>
<input>
<ID>IN_0</ID>597 </input>
<input>
<ID>IN_1</ID>604 </input>
<input>
<ID>IN_2</ID>605 </input>
<input>
<ID>IN_3</ID>546 </input>
<input>
<ID>IN_4</ID>598 </input>
<input>
<ID>IN_5</ID>608 </input>
<input>
<ID>IN_6</ID>609 </input>
<input>
<ID>IN_7</ID>610 </input>
<output>
<ID>OUT</ID>611 </output>
<input>
<ID>SEL_0</ID>599 </input>
<input>
<ID>SEL_1</ID>600 </input>
<input>
<ID>SEL_2</ID>601 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>695</ID>
<type>AA_AND2</type>
<position>124.5,-64.5</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>602 </input>
<output>
<ID>OUT</ID>597 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>696</ID>
<type>AE_SMALL_INVERTER</type>
<position>167,-0.5</position>
<input>
<ID>IN_0</ID>637 </input>
<output>
<ID>OUT_0</ID>628 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>697</ID>
<type>AE_SMALL_INVERTER</type>
<position>124.5,-55</position>
<input>
<ID>IN_0</ID>607 </input>
<output>
<ID>OUT_0</ID>598 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>698</ID>
<type>DA_FROM</type>
<position>117,-61</position>
<input>
<ID>IN_0</ID>604 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum11</lparam></gate>
<gate>
<ID>699</ID>
<type>AE_SMALL_INVERTER</type>
<position>166.5,23.5</position>
<input>
<ID>IN_0</ID>622 </input>
<output>
<ID>OUT_0</ID>613 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>700</ID>
<type>DA_FROM</type>
<position>117,-59</position>
<input>
<ID>IN_0</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr11</lparam></gate>
<gate>
<ID>701</ID>
<type>DA_FROM</type>
<position>117,-51</position>
<input>
<ID>IN_0</ID>609 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>702</ID>
<type>DA_FROM</type>
<position>117,-53</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>703</ID>
<type>DE_TO</type>
<position>-25,26</position>
<input>
<ID>IN_0</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr9</lparam></gate>
<gate>
<ID>705</ID>
<type>DA_FROM</type>
<position>117,-55</position>
<input>
<ID>IN_0</ID>607 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>706</ID>
<type>DA_FROM</type>
<position>117,-63</position>
<input>
<ID>IN_0</ID>603 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>707</ID>
<type>AI_MUX_8x1</type>
<position>178.5,-29.5</position>
<input>
<ID>IN_0</ID>642 </input>
<input>
<ID>IN_1</ID>649 </input>
<input>
<ID>IN_2</ID>650 </input>
<input>
<ID>IN_3</ID>591 </input>
<input>
<ID>IN_4</ID>643 </input>
<input>
<ID>IN_5</ID>660 </input>
<input>
<ID>IN_6</ID>661 </input>
<input>
<ID>IN_7</ID>662 </input>
<output>
<ID>OUT</ID>663 </output>
<input>
<ID>SEL_0</ID>644 </input>
<input>
<ID>SEL_1</ID>645 </input>
<input>
<ID>SEL_2</ID>646 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>709</ID>
<type>DA_FROM</type>
<position>136,-45.5</position>
<input>
<ID>IN_0</ID>600 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>710</ID>
<type>FF_GND</type>
<position>171,26</position>
<output>
<ID>OUT_0</ID>625 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>711</ID>
<type>FF_GND</type>
<position>171.5,2</position>
<output>
<ID>OUT_0</ID>640 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>713</ID>
<type>DA_FROM</type>
<position>159.5,-6.5</position>
<input>
<ID>IN_0</ID>634 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum13</lparam></gate>
<gate>
<ID>714</ID>
<type>DA_FROM</type>
<position>159.5,3.5</position>
<input>
<ID>IN_0</ID>639 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>715</ID>
<type>AA_AND2</type>
<position>166.5,14</position>
<input>
<ID>IN_0</ID>618 </input>
<input>
<ID>IN_1</ID>617 </input>
<output>
<ID>OUT</ID>612 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>717</ID>
<type>AE_SMALL_INVERTER</type>
<position>167,-28.5</position>
<input>
<ID>IN_0</ID>659 </input>
<output>
<ID>OUT_0</ID>643 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>718</ID>
<type>DA_FROM</type>
<position>159.5,-32.5</position>
<input>
<ID>IN_0</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr14</lparam></gate>
<gate>
<ID>719</ID>
<type>DA_FROM</type>
<position>159.5,-26.5</position>
<input>
<ID>IN_0</ID>660 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>720</ID>
<type>DA_FROM</type>
<position>159.5,-28.5</position>
<input>
<ID>IN_0</ID>659 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>721</ID>
<type>DA_FROM</type>
<position>159.5,-38.5</position>
<input>
<ID>IN_0</ID>647 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr14</lparam></gate>
<gate>
<ID>722</ID>
<type>DA_FROM</type>
<position>178.5,-19</position>
<input>
<ID>IN_0</ID>645 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>723</ID>
<type>DA_FROM</type>
<position>159,23.5</position>
<input>
<ID>IN_0</ID>622 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>724</ID>
<type>DA_FROM</type>
<position>159,13.5</position>
<input>
<ID>IN_0</ID>617 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr12</lparam></gate>
<gate>
<ID>725</ID>
<type>DA_FROM</type>
<position>178,33</position>
<input>
<ID>IN_0</ID>615 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>726</ID>
<type>AA_AND2</type>
<position>167,-10</position>
<input>
<ID>IN_0</ID>633 </input>
<input>
<ID>IN_1</ID>632 </input>
<output>
<ID>OUT</ID>627 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>727</ID>
<type>DA_FROM</type>
<position>159.5,-8.5</position>
<input>
<ID>IN_0</ID>633 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>728</ID>
<type>DA_FROM</type>
<position>178.5,9</position>
<input>
<ID>IN_0</ID>630 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>729</ID>
<type>DE_TO</type>
<position>183.5,-29.5</position>
<input>
<ID>IN_0</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin14</lparam></gate>
<gate>
<ID>730</ID>
<type>DA_FROM</type>
<position>159.5,-34.5</position>
<input>
<ID>IN_0</ID>649 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum14</lparam></gate>
<gate>
<ID>731</ID>
<type>DA_FROM</type>
<position>180.5,-19</position>
<input>
<ID>IN_0</ID>644 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>732</ID>
<type>FF_GND</type>
<position>172.5,-53</position>
<output>
<ID>OUT_0</ID>676 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>733</ID>
<type>AI_MUX_8x1</type>
<position>179.5,-56.5</position>
<input>
<ID>IN_0</ID>664 </input>
<input>
<ID>IN_1</ID>671 </input>
<input>
<ID>IN_2</ID>672 </input>
<input>
<ID>IN_3</ID>606 </input>
<input>
<ID>IN_4</ID>665 </input>
<input>
<ID>IN_5</ID>674 </input>
<input>
<ID>IN_6</ID>675 </input>
<input>
<ID>IN_7</ID>676 </input>
<output>
<ID>OUT</ID>677 </output>
<input>
<ID>SEL_0</ID>666 </input>
<input>
<ID>SEL_1</ID>667 </input>
<input>
<ID>SEL_2</ID>668 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>734</ID>
<type>AE_SMALL_INVERTER</type>
<position>168,-55.5</position>
<input>
<ID>IN_0</ID>673 </input>
<output>
<ID>OUT_0</ID>665 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>735</ID>
<type>DA_FROM</type>
<position>160.5,-59.5</position>
<input>
<ID>IN_0</ID>672 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr15</lparam></gate>
<gate>
<ID>736</ID>
<type>DA_FROM</type>
<position>160.5,-53.5</position>
<input>
<ID>IN_0</ID>674 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>737</ID>
<type>DA_FROM</type>
<position>160.5,-55.5</position>
<input>
<ID>IN_0</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>738</ID>
<type>DA_FROM</type>
<position>160.5,-65.5</position>
<input>
<ID>IN_0</ID>669 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr15</lparam></gate>
<gate>
<ID>739</ID>
<type>DA_FROM</type>
<position>181.5,-46</position>
<input>
<ID>IN_0</ID>666 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>772</ID>
<type>DE_TO</type>
<position>-58.5,-58.5</position>
<input>
<ID>IN_0</ID>716 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum10</lparam></gate>
<gate>
<ID>740</ID>
<type>DA_FROM</type>
<position>179.5,-46</position>
<input>
<ID>IN_0</ID>667 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>741</ID>
<type>DA_FROM</type>
<position>177.5,-46</position>
<input>
<ID>IN_0</ID>668 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>742</ID>
<type>DA_FROM</type>
<position>-13,-38</position>
<input>
<ID>IN_0</ID>705 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>743</ID>
<type>DA_FROM</type>
<position>-3.5,-38</position>
<input>
<ID>IN_0</ID>709 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr0</lparam></gate>
<gate>
<ID>744</ID>
<type>DA_FROM</type>
<position>-5.5,-38</position>
<input>
<ID>IN_0</ID>708 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr1</lparam></gate>
<gate>
<ID>745</ID>
<type>DA_FROM</type>
<position>-7.5,-38</position>
<input>
<ID>IN_0</ID>707 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr2</lparam></gate>
<gate>
<ID>770</ID>
<type>DE_TO</type>
<position>-35,-58.5</position>
<input>
<ID>IN_0</ID>720 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum6</lparam></gate>
<gate>
<ID>746</ID>
<type>DA_FROM</type>
<position>-9.5,-38</position>
<input>
<ID>IN_0</ID>706 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr3</lparam></gate>
<gate>
<ID>747</ID>
<type>DA_FROM</type>
<position>-25,-38</position>
<input>
<ID>IN_0</ID>701 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr4</lparam></gate>
<gate>
<ID>780</ID>
<type>DE_TO</type>
<position>-25,13</position>
<input>
<ID>IN_0</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr4</lparam></gate>
<gate>
<ID>748</ID>
<type>DA_FROM</type>
<position>-27,-38</position>
<input>
<ID>IN_0</ID>700 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr5</lparam></gate>
<gate>
<ID>749</ID>
<type>DA_FROM</type>
<position>-29,-38</position>
<input>
<ID>IN_0</ID>699 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr6</lparam></gate>
<gate>
<ID>774</ID>
<type>DE_TO</type>
<position>-82,-58.5</position>
<input>
<ID>IN_0</ID>714 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum14</lparam></gate>
<gate>
<ID>750</ID>
<type>DA_FROM</type>
<position>-31,-38</position>
<input>
<ID>IN_0</ID>698 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr7</lparam></gate>
<gate>
<ID>751</ID>
<type>DA_FROM</type>
<position>-49,-38</position>
<input>
<ID>IN_0</ID>693 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr8</lparam></gate>
<gate>
<ID>768</ID>
<type>DE_TO</type>
<position>-12.5,-58</position>
<input>
<ID>IN_0</ID>724 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum2</lparam></gate>
<gate>
<ID>752</ID>
<type>DA_FROM</type>
<position>-51,-38</position>
<input>
<ID>IN_0</ID>692 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr9</lparam></gate>
<gate>
<ID>753</ID>
<type>DA_FROM</type>
<position>-53,-38</position>
<input>
<ID>IN_0</ID>691 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr10</lparam></gate>
<gate>
<ID>778</ID>
<type>DE_TO</type>
<position>-25,7</position>
<input>
<ID>IN_0</ID>733 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr1</lparam></gate>
<gate>
<ID>754</ID>
<type>DA_FROM</type>
<position>-55,-38</position>
<input>
<ID>IN_0</ID>690 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr11</lparam></gate>
<gate>
<ID>755</ID>
<type>DA_FROM</type>
<position>-72.5,-38.5</position>
<input>
<ID>IN_0</ID>685 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr12</lparam></gate>
<gate>
<ID>788</ID>
<type>DA_FROM</type>
<position>71.5,-2</position>
<input>
<ID>IN_0</ID>456 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr5</lparam></gate>
<gate>
<ID>756</ID>
<type>DA_FROM</type>
<position>-74.5,-38.5</position>
<input>
<ID>IN_0</ID>684 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr13</lparam></gate>
<gate>
<ID>757</ID>
<type>DA_FROM</type>
<position>-76.5,-38.5</position>
<input>
<ID>IN_0</ID>683 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr14</lparam></gate>
<gate>
<ID>782</ID>
<type>DE_TO</type>
<position>-25,17</position>
<input>
<ID>IN_0</ID>728 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr6</lparam></gate>
<gate>
<ID>758</ID>
<type>DA_FROM</type>
<position>-78.5,-38.5</position>
<input>
<ID>IN_0</ID>682 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID dr15</lparam></gate>
<gate>
<ID>759</ID>
<type>DA_FROM</type>
<position>-15,-38</position>
<input>
<ID>IN_0</ID>704 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>776</ID>
<type>DE_TO</type>
<position>-25,11</position>
<input>
<ID>IN_0</ID>731 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr3</lparam></gate>
<gate>
<ID>760</ID>
<type>DA_FROM</type>
<position>-17,-38</position>
<input>
<ID>IN_0</ID>703 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>761</ID>
<type>DA_FROM</type>
<position>-34.5,-38</position>
<input>
<ID>IN_0</ID>697 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>786</ID>
<type>DA_FROM</type>
<position>25,-57</position>
<input>
<ID>IN_0</ID>432 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr3</lparam></gate>
<gate>
<ID>762</ID>
<type>DA_FROM</type>
<position>-38.5,-38</position>
<input>
<ID>IN_0</ID>695 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>763</ID>
<type>DA_FROM</type>
<position>-40.5,-38</position>
<input>
<ID>IN_0</ID>694 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>796</ID>
<type>DA_FROM</type>
<position>159.5,-2.5</position>
<input>
<ID>IN_0</ID>576 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr13</lparam></gate>
<gate>
<ID>764</ID>
<type>DA_FROM</type>
<position>-59,-38</position>
<input>
<ID>IN_0</ID>688 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>765</ID>
<type>DA_FROM</type>
<position>-63,-38</position>
<input>
<ID>IN_0</ID>687 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>790</ID>
<type>DA_FROM</type>
<position>72.5,-57</position>
<input>
<ID>IN_0</ID>486 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr7</lparam></gate>
<gate>
<ID>766</ID>
<type>DA_FROM</type>
<position>-81.5,-38.5</position>
<input>
<ID>IN_0</ID>678 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>767</ID>
<type>DA_FROM</type>
<position>-85.5,-38.5</position>
<input>
<ID>IN_0</ID>680 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>784</ID>
<type>DA_FROM</type>
<position>24,-2</position>
<input>
<ID>IN_0</ID>414 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr1</lparam></gate>
<gate>
<ID>769</ID>
<type>DE_TO</type>
<position>-31,-58.5</position>
<input>
<ID>IN_0</ID>722 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum4</lparam></gate>
<gate>
<ID>771</ID>
<type>DE_TO</type>
<position>-54.5,-58.5</position>
<input>
<ID>IN_0</ID>718 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum8</lparam></gate>
<gate>
<ID>773</ID>
<type>DE_TO</type>
<position>-78,-58.5</position>
<input>
<ID>IN_0</ID>711 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum12</lparam></gate>
<gate>
<ID>775</ID>
<type>DA_FROM</type>
<position>-45,4.5</position>
<input>
<ID>IN_0</ID>735 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>777</ID>
<type>DE_TO</type>
<position>-25,5</position>
<input>
<ID>IN_0</ID>734 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr0</lparam></gate>
<gate>
<ID>779</ID>
<type>DE_TO</type>
<position>-25,9</position>
<input>
<ID>IN_0</ID>732 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr2</lparam></gate>
<gate>
<ID>781</ID>
<type>DE_TO</type>
<position>-25,15</position>
<input>
<ID>IN_0</ID>729 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr5</lparam></gate>
<gate>
<ID>783</ID>
<type>DE_TO</type>
<position>-25,19</position>
<input>
<ID>IN_0</ID>727 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr7</lparam></gate>
<gate>
<ID>785</ID>
<type>DA_FROM</type>
<position>24,-30</position>
<input>
<ID>IN_0</ID>415 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr2</lparam></gate>
<gate>
<ID>787</ID>
<type>DA_FROM</type>
<position>71,22</position>
<input>
<ID>IN_0</ID>433 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr4</lparam></gate>
<gate>
<ID>789</ID>
<type>DA_FROM</type>
<position>71.5,-30</position>
<input>
<ID>IN_0</ID>471 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr6</lparam></gate>
<gate>
<ID>791</ID>
<type>DA_FROM</type>
<position>115.5,22</position>
<input>
<ID>IN_0</ID>501 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr8</lparam></gate>
<gate>
<ID>795</ID>
<type>DA_FROM</type>
<position>159,21.5</position>
<input>
<ID>IN_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr12</lparam></gate>
<gate>
<ID>797</ID>
<type>DA_FROM</type>
<position>159.5,-30.5</position>
<input>
<ID>IN_0</ID>591 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr14</lparam></gate>
<gate>
<ID>799</ID>
<type>DE_TO</type>
<position>-93.5,-49</position>
<input>
<ID>IN_0</ID>621 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Cout</lparam></gate>
<gate>
<ID>803</ID>
<type>BV_4x1_BUS_END</type>
<position>-50,14</position>
<input>
<ID>IN_0</ID>402 </input>
<input>
<ID>IN_1</ID>403 </input>
<input>
<ID>IN_2</ID>404 </input>
<input>
<ID>IN_3</ID>405 </input>
<input>
<ID>OUT</ID>746 747 748 749 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>807</ID>
<type>DE_TO</type>
<position>-25,34</position>
<input>
<ID>IN_0</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr13</lparam></gate>
<gate>
<ID>811</ID>
<type>BV_4x1_BUS_END</type>
<position>-50,18</position>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>815</ID>
<type>FF_GND</type>
<position>-29,22</position>
<output>
<ID>OUT_0</ID>397 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>621 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-91.5,-49,-89,-49</points>
<connection>
<GID>486</GID>
<name>carry_out</name></connection>
<connection>
<GID>799</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>444 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,25.5,33,28</points>
<intersection>25.5 2</intersection>
<intersection>28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,28,33,28</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,25.5,39.5,25.5</points>
<connection>
<GID>483</GID>
<name>IN_6</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>557 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,13.5,118.5,14</points>
<intersection>13.5 1</intersection>
<intersection>14 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118.5,13.5,120,13.5</points>
<connection>
<GID>639</GID>
<name>IN_1</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>117.5,14,118.5,14</points>
<connection>
<GID>664</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>476 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-29,46,-29</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<connection>
<GID>489</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>413 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,13.5,-40,13.5</points>
<connection>
<GID>804</GID>
<name>OUT_5</name></connection>
<connection>
<GID>816</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>405 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48,15.5,-48,15.5</points>
<connection>
<GID>804</GID>
<name>IN_7</name></connection>
<connection>
<GID>803</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>740 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75,5.5,-75,7</points>
<intersection>5.5 1</intersection>
<intersection>7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76,5.5,-75,5.5</points>
<connection>
<GID>801</GID>
<name>OUT_0</name></connection>
<intersection>-75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-75,7,-73.5,7</points>
<connection>
<GID>802</GID>
<name>IN_0</name></connection>
<intersection>-75 0</intersection></hsegment></shape></wire>
<wire>
<ID>746 747 748 749 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,8.5,-62,14</points>
<intersection>8.5 1</intersection>
<intersection>14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69.5,8.5,-62,8.5</points>
<connection>
<GID>802</GID>
<name>OUT</name></connection>
<intersection>-62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-62,14,-52,14</points>
<connection>
<GID>803</GID>
<name>OUT</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>455 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-4,33,-2.5</points>
<intersection>-4 1</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-4,33,-4</points>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-2.5,40,-2.5</points>
<connection>
<GID>473</GID>
<name>IN_2</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>546 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-57,126,-56.5</points>
<intersection>-57 2</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,-56.5,133,-56.5</points>
<connection>
<GID>694</GID>
<name>IN_3</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119,-57,126,-57</points>
<connection>
<GID>794</GID>
<name>IN_0</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>738 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75,7.5,-75,8</points>
<intersection>7.5 1</intersection>
<intersection>8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76,7.5,-75,7.5</points>
<connection>
<GID>801</GID>
<name>OUT_1</name></connection>
<intersection>-75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-75,8,-73.5,8</points>
<connection>
<GID>802</GID>
<name>IN_1</name></connection>
<intersection>-75 0</intersection></hsegment></shape></wire>
<wire>
<ID>739 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75,9,-75,9.5</points>
<intersection>9 2</intersection>
<intersection>9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76,9.5,-75,9.5</points>
<connection>
<GID>801</GID>
<name>OUT_2</name></connection>
<intersection>-75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-75,9,-73.5,9</points>
<connection>
<GID>802</GID>
<name>IN_2</name></connection>
<intersection>-75 0</intersection></hsegment></shape></wire>
<wire>
<ID>737 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75,10,-75,11.5</points>
<intersection>10 2</intersection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76,11.5,-75,11.5</points>
<connection>
<GID>801</GID>
<name>OUT_3</name></connection>
<intersection>-75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-75,10,-73.5,10</points>
<connection>
<GID>802</GID>
<name>IN_3</name></connection>
<intersection>-75 0</intersection></hsegment></shape></wire>
<wire>
<ID>623 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,24,168,25.5</points>
<intersection>24 1</intersection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,24,175,24</points>
<connection>
<GID>678</GID>
<name>IN_5</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161,25.5,168,25.5</points>
<connection>
<GID>540</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment></shape></wire>
<wire>
<ID>458 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,0.5,33,2</points>
<intersection>0.5 1</intersection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,0.5,40,0.5</points>
<connection>
<GID>473</GID>
<name>IN_5</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,2,33,2</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>559 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,18,126,20.5</points>
<intersection>18 2</intersection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,20.5,131.5,20.5</points>
<connection>
<GID>637</GID>
<name>IN_1</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>117.5,18,126,18</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>583 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-28.5,128.5,-28</points>
<intersection>-28.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128.5,-28.5,132,-28.5</points>
<connection>
<GID>643</GID>
<name>IN_4</name></connection>
<intersection>128.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125.5,-28,128.5,-28</points>
<connection>
<GID>645</GID>
<name>OUT_0</name></connection>
<intersection>128.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>418 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32,-16.5,-32,-13.5</points>
<intersection>-16.5 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32,-16.5,-23,-16.5</points>
<connection>
<GID>504</GID>
<name>IN_5</name></connection>
<intersection>-32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-36.5,-13.5,-32,-13.5</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<intersection>-32 0</intersection></hsegment></shape></wire>
<wire>
<ID>613 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171.5,23,171.5,23.5</points>
<intersection>23 1</intersection>
<intersection>23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171.5,23,175,23</points>
<connection>
<GID>678</GID>
<name>IN_4</name></connection>
<intersection>171.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>168.5,23.5,171.5,23.5</points>
<connection>
<GID>699</GID>
<name>OUT_0</name></connection>
<intersection>171.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>436 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,28.5,40.5,31.5</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<intersection>28.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>40.5,28.5,41.5,28.5</points>
<connection>
<GID>483</GID>
<name>SEL_2</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>558 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>117.5,16,120,16</points>
<connection>
<GID>662</GID>
<name>IN_0</name></connection>
<intersection>120 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>120,15.5,120,16</points>
<connection>
<GID>639</GID>
<name>IN_0</name></connection>
<intersection>16 1</intersection></vsegment></shape></wire>
<wire>
<ID>451 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,4.5,41,7.5</points>
<connection>
<GID>520</GID>
<name>IN_0</name></connection>
<intersection>4.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>41,4.5,42,4.5</points>
<connection>
<GID>473</GID>
<name>SEL_2</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>686 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62.5,-46,-62.5,-43</points>
<connection>
<GID>507</GID>
<name>IN_3</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-65,-43,-62.5,-43</points>
<intersection>-65 3</intersection>
<intersection>-62.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-65,-43,-65,-40</points>
<connection>
<GID>641</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>445 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,26.5,35.5,27.5</points>
<connection>
<GID>464</GID>
<name>OUT_0</name></connection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,26.5,39.5,26.5</points>
<connection>
<GID>483</GID>
<name>IN_7</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>571 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,4.5,133,7.5</points>
<connection>
<GID>677</GID>
<name>IN_0</name></connection>
<intersection>4.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>133,4.5,134,4.5</points>
<connection>
<GID>630</GID>
<name>SEL_2</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>422 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-21.5,-30,-20.5</points>
<intersection>-21.5 1</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-21.5,-30,-21.5</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-30,-20.5,-23,-20.5</points>
<connection>
<GID>504</GID>
<name>IN_1</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>641 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-1.5,181.5,-1.5</points>
<connection>
<GID>681</GID>
<name>IN_0</name></connection>
<connection>
<GID>712</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>464 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-23.5,44,-22</points>
<connection>
<GID>489</GID>
<name>SEL_0</name></connection>
<intersection>-22 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>45,-22,45,-20.5</points>
<connection>
<GID>526</GID>
<name>IN_0</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>44,-22,45,-22</points>
<intersection>44 0</intersection>
<intersection>45 1</intersection></hsegment></shape></wire>
<wire>
<ID>400 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48,11.5,-48,11.5</points>
<connection>
<GID>685</GID>
<name>IN_3</name></connection>
<connection>
<GID>804</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>577 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118,0,121.5,0</points>
<connection>
<GID>671</GID>
<name>IN_0</name></connection>
<connection>
<GID>631</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>425 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17,-19,-10.5,-19</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>-17 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-17,-19.5,-17,-19</points>
<connection>
<GID>504</GID>
<name>OUT_2</name></connection>
<intersection>-19 1</intersection></vsegment></shape></wire>
<wire>
<ID>568 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-0.5,128.5,0</points>
<intersection>-0.5 1</intersection>
<intersection>0 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128.5,-0.5,132,-0.5</points>
<connection>
<GID>630</GID>
<name>IN_4</name></connection>
<intersection>128.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125.5,0,128.5,0</points>
<connection>
<GID>631</GID>
<name>OUT_0</name></connection>
<intersection>128.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>421 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36.5,-19.5,-23,-19.5</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<connection>
<GID>504</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>461 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-1,46,-1</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<connection>
<GID>473</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>732 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,9,-28,10.5</points>
<intersection>9 1</intersection>
<intersection>10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-28,9,-27,9</points>
<connection>
<GID>779</GID>
<name>IN_0</name></connection>
<intersection>-28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,10.5,-28,10.5</points>
<connection>
<GID>817</GID>
<name>IN_2</name></connection>
<intersection>-28 0</intersection></hsegment></shape></wire>
<wire>
<ID>397 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,23,-29,38</points>
<connection>
<GID>815</GID>
<name>OUT_0</name></connection>
<intersection>24 16</intersection>
<intersection>26 15</intersection>
<intersection>28 14</intersection>
<intersection>30 13</intersection>
<intersection>32 12</intersection>
<intersection>34 11</intersection>
<intersection>36 10</intersection>
<intersection>38 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-29,38,-27,38</points>
<connection>
<GID>805</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-29,36,-27,36</points>
<connection>
<GID>806</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-29,34,-27,34</points>
<connection>
<GID>807</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-29,32,-27,32</points>
<connection>
<GID>580</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-29,30,-27,30</points>
<connection>
<GID>808</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-29,28,-27,28</points>
<connection>
<GID>809</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-29,26,-27,26</points>
<connection>
<GID>703</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-29,24,-27,24</points>
<connection>
<GID>810</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>510 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,4.5,90.5,7.5</points>
<connection>
<GID>550</GID>
<name>SEL_1</name></connection>
<connection>
<GID>598</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>531 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-30,125,-29.5</points>
<intersection>-30 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-29.5,132,-29.5</points>
<connection>
<GID>643</GID>
<name>IN_3</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>118,-30,125,-30</points>
<connection>
<GID>793</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>446 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,23,45.5,23</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<connection>
<GID>483</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>453 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-8.5,27,-8</points>
<intersection>-8.5 2</intersection>
<intersection>-8 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27,-8.5,28.5,-8.5</points>
<connection>
<GID>514</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26,-8,27,-8</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>435 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,28.5,42.5,31.5</points>
<connection>
<GID>483</GID>
<name>SEL_1</name></connection>
<connection>
<GID>512</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>606 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-57.5,169.5,-57</points>
<intersection>-57.5 2</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-57,176.5,-57</points>
<connection>
<GID>733</GID>
<name>IN_3</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-57.5,169.5,-57.5</points>
<connection>
<GID>798</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>449 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,4.5,44,6</points>
<connection>
<GID>473</GID>
<name>SEL_0</name></connection>
<intersection>6 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>45,6,45,7.5</points>
<connection>
<GID>518</GID>
<name>IN_0</name></connection>
<intersection>6 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>44,6,45,6</points>
<intersection>44 0</intersection>
<intersection>45 1</intersection></hsegment></shape></wire>
<wire>
<ID>592 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118,-28,121.5,-28</points>
<connection>
<GID>654</GID>
<name>IN_0</name></connection>
<connection>
<GID>645</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>597 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,-64.5,132.5,-59.5</points>
<intersection>-64.5 2</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-59.5,133,-59.5</points>
<connection>
<GID>694</GID>
<name>IN_0</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-64.5,132.5,-64.5</points>
<connection>
<GID>695</GID>
<name>OUT</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>420 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34.5,-18.5,-34.5,-17.5</points>
<intersection>-18.5 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-18.5,-23,-18.5</points>
<connection>
<GID>504</GID>
<name>IN_3</name></connection>
<intersection>-34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-36.5,-17.5,-34.5,-17.5</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>-34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>460 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,2.5,36,3.5</points>
<connection>
<GID>469</GID>
<name>OUT_0</name></connection>
<intersection>2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,2.5,40,2.5</points>
<connection>
<GID>473</GID>
<name>IN_7</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>603 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-63.5,120,-63</points>
<intersection>-63.5 2</intersection>
<intersection>-63 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>120,-63.5,121.5,-63.5</points>
<connection>
<GID>695</GID>
<name>IN_0</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>119,-63,120,-63</points>
<connection>
<GID>706</GID>
<name>IN_0</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>454 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-6,34.5,-3.5</points>
<intersection>-6 2</intersection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-3.5,40,-3.5</points>
<connection>
<GID>473</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-6,34.5,-6</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>539 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-50.5,92.5,-49</points>
<connection>
<GID>609</GID>
<name>SEL_0</name></connection>
<intersection>-49 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>93.5,-49,93.5,-47.5</points>
<connection>
<GID>619</GID>
<name>IN_0</name></connection>
<intersection>-49 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-49,93.5,-49</points>
<intersection>92.5 0</intersection>
<intersection>93.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>419 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-17.5,-33.5,-15.5</points>
<intersection>-17.5 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-15.5,-33.5,-15.5</points>
<connection>
<GID>470</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33.5,-17.5,-23,-17.5</points>
<connection>
<GID>504</GID>
<name>IN_4</name></connection>
<intersection>-33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>447 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-9.5,39.5,-4.5</points>
<intersection>-9.5 2</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-4.5,40,-4.5</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-9.5,39.5,-9.5</points>
<connection>
<GID>514</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>563 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,24.5,124.5,26</points>
<intersection>24.5 1</intersection>
<intersection>26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,24.5,131.5,24.5</points>
<connection>
<GID>637</GID>
<name>IN_5</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>117.5,26,124.5,26</points>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>414 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-2,33,-1.5</points>
<intersection>-2 2</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-1.5,40,-1.5</points>
<connection>
<GID>473</GID>
<name>IN_3</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-2,33,-2</points>
<connection>
<GID>784</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>448 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-0.5,36.5,0</points>
<intersection>-0.5 1</intersection>
<intersection>0 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-0.5,40,-0.5</points>
<connection>
<GID>473</GID>
<name>IN_4</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,0,36.5,0</points>
<connection>
<GID>475</GID>
<name>OUT_0</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>459 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,1.5,33.5,4</points>
<intersection>1.5 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,4,33.5,4</points>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,1.5,40,1.5</points>
<connection>
<GID>473</GID>
<name>IN_6</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>615 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178,28,178,31</points>
<connection>
<GID>678</GID>
<name>SEL_1</name></connection>
<connection>
<GID>725</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>450 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,4.5,43,7.5</points>
<connection>
<GID>473</GID>
<name>SEL_1</name></connection>
<connection>
<GID>519</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>552 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,14.5,131,19.5</points>
<intersection>14.5 2</intersection>
<intersection>19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,19.5,131.5,19.5</points>
<connection>
<GID>637</GID>
<name>IN_0</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>126,14.5,131,14.5</points>
<connection>
<GID>639</GID>
<name>OUT</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>417 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-15.5,-30,-11.5</points>
<intersection>-15.5 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-11.5,-30,-11.5</points>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-30,-15.5,-23,-15.5</points>
<connection>
<GID>504</GID>
<name>IN_6</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>401 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48,9.5,-48,9.5</points>
<connection>
<GID>685</GID>
<name>IN_1</name></connection>
<connection>
<GID>804</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>736 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,17.5,-44,21.5</points>
<connection>
<GID>804</GID>
<name>count_enable</name></connection>
<intersection>21.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-44,21.5,-39.5,21.5</points>
<connection>
<GID>813</GID>
<name>OUT_0</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>457 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,0,29.5,0</points>
<connection>
<GID>516</GID>
<name>IN_0</name></connection>
<connection>
<GID>475</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>645 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-24,178.5,-21</points>
<connection>
<GID>707</GID>
<name>SEL_1</name></connection>
<connection>
<GID>722</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>468 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-36.5,27,-36</points>
<intersection>-36.5 2</intersection>
<intersection>-36 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27,-36.5,28.5,-36.5</points>
<connection>
<GID>522</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26,-36,27,-36</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>427 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-23,-14,-21.5</points>
<intersection>-23 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17,-21.5,-14,-21.5</points>
<connection>
<GID>504</GID>
<name>OUT_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-14,-23,-10.5,-23</points>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>726 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-55,-10,-54</points>
<connection>
<GID>490</GID>
<name>OUT_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-8.5,-56,-8.5,-55</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-10,-55,-8.5,-55</points>
<intersection>-10 0</intersection>
<intersection>-8.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>580 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,2.5,128,3.5</points>
<connection>
<GID>627</GID>
<name>OUT_0</name></connection>
<intersection>2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,2.5,132,2.5</points>
<connection>
<GID>630</GID>
<name>IN_7</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>426 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-21,-14,-20.5</points>
<intersection>-21 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17,-20.5,-14,-20.5</points>
<connection>
<GID>504</GID>
<name>OUT_1</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-14,-21,-10.5,-21</points>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>587 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-38.5,119,-38</points>
<intersection>-38.5 1</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-38.5,120.5,-38.5</points>
<connection>
<GID>680</GID>
<name>IN_1</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>118,-38,119,-38</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>423 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-23.5,-29,-21.5</points>
<intersection>-23.5 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29,-21.5,-23,-21.5</points>
<connection>
<GID>504</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-36.5,-23.5,-29,-23.5</points>
<connection>
<GID>482</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>585 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-23.5,135,-20.5</points>
<connection>
<GID>643</GID>
<name>SEL_1</name></connection>
<connection>
<GID>659</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>408 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,14.5,39,19.5</points>
<intersection>14.5 2</intersection>
<intersection>19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,19.5,39.5,19.5</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,14.5,39,14.5</points>
<connection>
<GID>484</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>439 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,18,34,20.5</points>
<intersection>18 2</intersection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,20.5,39.5,20.5</points>
<connection>
<GID>483</GID>
<name>IN_1</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,18,34,18</points>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>617 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,13,162,13.5</points>
<intersection>13 1</intersection>
<intersection>13.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162,13,163.5,13</points>
<connection>
<GID>715</GID>
<name>IN_1</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>161,13.5,162,13.5</points>
<connection>
<GID>724</GID>
<name>IN_0</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>440 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,20,32.5,21.5</points>
<intersection>20 1</intersection>
<intersection>21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,20,32.5,20</points>
<connection>
<GID>496</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,21.5,39.5,21.5</points>
<connection>
<GID>483</GID>
<name>IN_2</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>648 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162.5,-37,162.5,-36.5</points>
<intersection>-37 2</intersection>
<intersection>-36.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-37,164,-37</points>
<connection>
<GID>555</GID>
<name>IN_0</name></connection>
<intersection>162.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>161.5,-36.5,162.5,-36.5</points>
<connection>
<GID>584</GID>
<name>IN_0</name></connection>
<intersection>162.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>441 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,22,32.5,22.5</points>
<intersection>22 2</intersection>
<intersection>22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,22.5,39.5,22.5</points>
<connection>
<GID>483</GID>
<name>IN_3</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,22,32.5,22</points>
<connection>
<GID>502</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>431 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,23.5,36,24</points>
<intersection>23.5 1</intersection>
<intersection>24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,23.5,39.5,23.5</points>
<connection>
<GID>483</GID>
<name>IN_4</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,24,36,24</points>
<connection>
<GID>492</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>443 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,24.5,32.5,26</points>
<intersection>24.5 1</intersection>
<intersection>26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,24.5,39.5,24.5</points>
<connection>
<GID>483</GID>
<name>IN_5</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,26,32.5,26</points>
<connection>
<GID>500</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>434 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,28.5,43.5,30</points>
<connection>
<GID>483</GID>
<name>SEL_0</name></connection>
<intersection>30 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>44.5,30,44.5,31.5</points>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<intersection>30 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>43.5,30,44.5,30</points>
<intersection>43.5 0</intersection>
<intersection>44.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>745 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45,17.5,-45,22.5</points>
<connection>
<GID>804</GID>
<name>load</name></connection>
<connection>
<GID>814</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>562 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>117.5,24,121,24</points>
<connection>
<GID>661</GID>
<name>IN_0</name></connection>
<connection>
<GID>646</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>438 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,15.5,26.5,16</points>
<intersection>15.5 2</intersection>
<intersection>16 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>26.5,15.5,28,15.5</points>
<connection>
<GID>484</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25.5,16,26.5,16</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>644 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-24,179.5,-22.5</points>
<connection>
<GID>707</GID>
<name>SEL_0</name></connection>
<intersection>-22.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>180.5,-22.5,180.5,-21</points>
<connection>
<GID>731</GID>
<name>IN_0</name></connection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>179.5,-22.5,180.5,-22.5</points>
<intersection>179.5 0</intersection>
<intersection>180.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>437 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,13.5,26.5,14</points>
<intersection>13.5 1</intersection>
<intersection>14 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,13.5,28,13.5</points>
<connection>
<GID>484</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25.5,14,26.5,14</points>
<connection>
<GID>510</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>452 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-10.5,27,-10</points>
<intersection>-10.5 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-10.5,28.5,-10.5</points>
<connection>
<GID>514</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-10,27,-10</points>
<connection>
<GID>485</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>723 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-56,-14.5,-55</points>
<connection>
<GID>635</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-13,-55,-13,-54</points>
<connection>
<GID>490</GID>
<name>OUT_3</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-14.5,-55,-13,-55</points>
<intersection>-14.5 0</intersection>
<intersection>-13 1</intersection></hsegment></shape></wire>
<wire>
<ID>678 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-83,-46,-83,-43</points>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-81.5,-43,-81.5,-40.5</points>
<connection>
<GID>766</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-83,-43,-81.5,-43</points>
<intersection>-83 0</intersection>
<intersection>-81.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>679 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84,-46,-84,-43</points>
<connection>
<GID>486</GID>
<name>IN_1</name></connection>
<intersection>-43 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-83.5,-43,-83.5,-40.5</points>
<connection>
<GID>632</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-84,-43,-83.5,-43</points>
<intersection>-84 0</intersection>
<intersection>-83.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>680 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-85.5,-43,-85.5,-40.5</points>
<connection>
<GID>767</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-85,-46,-85,-43</points>
<connection>
<GID>486</GID>
<name>IN_2</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-85.5,-43,-85,-43</points>
<intersection>-85.5 0</intersection>
<intersection>-85 1</intersection></hsegment></shape></wire>
<wire>
<ID>504 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,25.5,80.5,28</points>
<intersection>25.5 2</intersection>
<intersection>28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,28,80.5,28</points>
<connection>
<GID>575</GID>
<name>IN_0</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80.5,25.5,87,25.5</points>
<connection>
<GID>557</GID>
<name>IN_6</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>681 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86,-46,-86,-43</points>
<connection>
<GID>486</GID>
<name>IN_3</name></connection>
<intersection>-43 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-87.5,-43,-87.5,-40.5</points>
<connection>
<GID>623</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-43,-86,-43</points>
<intersection>-87.5 1</intersection>
<intersection>-86 0</intersection></hsegment></shape></wire>
<wire>
<ID>508 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-0.5,84,0</points>
<intersection>-0.5 1</intersection>
<intersection>0 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-0.5,87.5,-0.5</points>
<connection>
<GID>550</GID>
<name>IN_4</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81,0,84,0</points>
<connection>
<GID>551</GID>
<name>OUT_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>685 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72.5,-43,-72.5,-40.5</points>
<connection>
<GID>755</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-73,-46,-73,-43</points>
<intersection>-46 3</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-73,-43,-72.5,-43</points>
<intersection>-73 1</intersection>
<intersection>-72.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-76,-46,-73,-46</points>
<connection>
<GID>486</GID>
<name>IN_B_0</name></connection>
<intersection>-73 1</intersection></hsegment></shape></wire>
<wire>
<ID>684 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77,-46,-77,-43</points>
<connection>
<GID>486</GID>
<name>IN_B_1</name></connection>
<intersection>-43 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-74.5,-43,-74.5,-40.5</points>
<connection>
<GID>756</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-77,-43,-74.5,-43</points>
<intersection>-77 0</intersection>
<intersection>-74.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>683 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,-43,-77.5,-40.5</points>
<intersection>-43 2</intersection>
<intersection>-40.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-78,-46,-78,-43</points>
<connection>
<GID>486</GID>
<name>IN_B_2</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-78,-43,-77.5,-43</points>
<intersection>-78 1</intersection>
<intersection>-77.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-77.5,-40.5,-76.5,-40.5</points>
<connection>
<GID>757</GID>
<name>IN_0</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>682 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78.5,-46,-78.5,-40.5</points>
<connection>
<GID>758</GID>
<name>IN_0</name></connection>
<intersection>-46 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-79,-46,-78.5,-46</points>
<connection>
<GID>486</GID>
<name>IN_B_3</name></connection>
<intersection>-78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>430 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-73,-49,-65.5,-49</points>
<connection>
<GID>486</GID>
<name>carry_in</name></connection>
<connection>
<GID>507</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>711 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,-56.5,-78,-55</points>
<connection>
<GID>773</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-79.5,-55,-79.5,-54</points>
<connection>
<GID>486</GID>
<name>OUT_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-79.5,-55,-78,-55</points>
<intersection>-79.5 1</intersection>
<intersection>-78 0</intersection></hsegment></shape></wire>
<wire>
<ID>505 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,26.5,83,27.5</points>
<connection>
<GID>544</GID>
<name>OUT_0</name></connection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,26.5,87,26.5</points>
<connection>
<GID>557</GID>
<name>IN_7</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>712 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80,-56.5,-80,-55</points>
<connection>
<GID>660</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-80.5,-55,-80.5,-54</points>
<connection>
<GID>486</GID>
<name>OUT_1</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-80.5,-55,-80,-55</points>
<intersection>-80.5 1</intersection>
<intersection>-80 0</intersection></hsegment></shape></wire>
<wire>
<ID>714 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-82,-56.5,-82,-55</points>
<connection>
<GID>774</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-81.5,-55,-81.5,-54</points>
<connection>
<GID>486</GID>
<name>OUT_2</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-82,-55,-81.5,-55</points>
<intersection>-82 0</intersection>
<intersection>-81.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>713 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84,-56.5,-84,-55</points>
<connection>
<GID>672</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-82.5,-55,-82.5,-54</points>
<connection>
<GID>486</GID>
<name>OUT_3</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-84,-55,-82.5,-55</points>
<intersection>-84 0</intersection>
<intersection>-82.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>475 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-25.5,36,-24.5</points>
<connection>
<GID>487</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-25.5,40,-25.5</points>
<connection>
<GID>489</GID>
<name>IN_7</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>554 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,28.5,135.5,30</points>
<connection>
<GID>637</GID>
<name>SEL_0</name></connection>
<intersection>30 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>136.5,30,136.5,31.5</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<intersection>30 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>135.5,30,136.5,30</points>
<intersection>135.5 0</intersection>
<intersection>136.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>697 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-46,-36,-43</points>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-36,-43,-34.5,-43</points>
<intersection>-36 0</intersection>
<intersection>-34.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-34.5,-43,-34.5,-40</points>
<connection>
<GID>761</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>696 </ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-37,-46,-37,-43</points>
<connection>
<GID>488</GID>
<name>IN_1</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-37,-43,-36.5,-43</points>
<intersection>-37 1</intersection>
<intersection>-36.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-36.5,-43,-36.5,-40</points>
<connection>
<GID>620</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>695 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38,-46,-38,-43</points>
<connection>
<GID>488</GID>
<name>IN_2</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-38.5,-43,-38,-43</points>
<intersection>-38.5 3</intersection>
<intersection>-38 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-38.5,-43,-38.5,-40</points>
<connection>
<GID>762</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>694 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39,-46,-39,-43</points>
<connection>
<GID>488</GID>
<name>IN_3</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-40.5,-43,-39,-43</points>
<intersection>-40.5 3</intersection>
<intersection>-39 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-40.5,-43,-40.5,-40</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>701 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-46,-29,-44.5</points>
<connection>
<GID>488</GID>
<name>IN_B_0</name></connection>
<intersection>-44.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-25,-44.5,-25,-40</points>
<connection>
<GID>747</GID>
<name>IN_0</name></connection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-29,-44.5,-25,-44.5</points>
<intersection>-29 0</intersection>
<intersection>-25 1</intersection></hsegment></shape></wire>
<wire>
<ID>700 </ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-30,-46,-30,-43</points>
<connection>
<GID>488</GID>
<name>IN_B_1</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-30,-43,-27,-43</points>
<intersection>-30 1</intersection>
<intersection>-27 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-27,-43,-27,-40</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>699 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,-46,-31,-43</points>
<connection>
<GID>488</GID>
<name>IN_B_2</name></connection>
<intersection>-43 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-30.5,-43,-30.5,-40</points>
<intersection>-43 2</intersection>
<intersection>-40 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-31,-43,-30.5,-43</points>
<intersection>-31 0</intersection>
<intersection>-30.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-30.5,-40,-29,-40</points>
<connection>
<GID>749</GID>
<name>IN_0</name></connection>
<intersection>-30.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>698 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32,-46,-32,-40</points>
<connection>
<GID>488</GID>
<name>IN_B_3</name></connection>
<intersection>-40 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-32,-40,-31,-40</points>
<connection>
<GID>750</GID>
<name>IN_0</name></connection>
<intersection>-32 0</intersection></hsegment></shape></wire>
<wire>
<ID>605 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-59,126,-57.5</points>
<intersection>-59 1</intersection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-59,126,-59</points>
<connection>
<GID>700</GID>
<name>IN_0</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>126,-57.5,133,-57.5</points>
<connection>
<GID>694</GID>
<name>IN_2</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>428 </ID>
<shape>
<hsegment>
<ID>15</ID>
<points>-26,-49,-19.5,-49</points>
<connection>
<GID>488</GID>
<name>carry_in</name></connection>
<connection>
<GID>490</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>722 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,-56.5,-31,-55</points>
<connection>
<GID>769</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-32.5,-55,-32.5,-54</points>
<connection>
<GID>488</GID>
<name>OUT_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-32.5,-55,-31,-55</points>
<intersection>-32.5 1</intersection>
<intersection>-31 0</intersection></hsegment></shape></wire>
<wire>
<ID>721 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-55,-33.5,-54</points>
<connection>
<GID>488</GID>
<name>OUT_1</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-33,-56.5,-33,-55</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-33.5,-55,-33,-55</points>
<intersection>-33.5 0</intersection>
<intersection>-33 1</intersection></hsegment></shape></wire>
<wire>
<ID>720 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-56.5,-35,-55</points>
<connection>
<GID>770</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-34.5,-55,-34.5,-54</points>
<connection>
<GID>488</GID>
<name>OUT_2</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-35,-55,-34.5,-55</points>
<intersection>-35 0</intersection>
<intersection>-34.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>719 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-55,-35.5,-54</points>
<connection>
<GID>488</GID>
<name>OUT_3</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-37,-56.5,-37,-55</points>
<connection>
<GID>663</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-37,-55,-35.5,-55</points>
<intersection>-37 1</intersection>
<intersection>-35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>429 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-49.5,-49,-42,-49</points>
<connection>
<GID>507</GID>
<name>carry_in</name></connection>
<connection>
<GID>488</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>611 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-56,139,-56</points>
<connection>
<GID>692</GID>
<name>IN_0</name></connection>
<connection>
<GID>694</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>462 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-37.5,39.5,-32.5</points>
<intersection>-37.5 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-32.5,40,-32.5</points>
<connection>
<GID>489</GID>
<name>IN_0</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-37.5,39.5,-37.5</points>
<connection>
<GID>522</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>469 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-34,34.5,-31.5</points>
<intersection>-34 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-31.5,40,-31.5</points>
<connection>
<GID>489</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-34,34.5,-34</points>
<connection>
<GID>523</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>619 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,17.5,169.5,20</points>
<intersection>17.5 2</intersection>
<intersection>20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,20,175,20</points>
<connection>
<GID>678</GID>
<name>IN_1</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161,17.5,169.5,17.5</points>
<connection>
<GID>690</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>470 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-32,33,-30.5</points>
<intersection>-32 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-32,33,-32</points>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-30.5,40,-30.5</points>
<connection>
<GID>489</GID>
<name>IN_2</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>415 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-30,33,-29.5</points>
<intersection>-30 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-29.5,40,-29.5</points>
<connection>
<GID>489</GID>
<name>IN_3</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-30,33,-30</points>
<connection>
<GID>785</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>463 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-28.5,36.5,-28</points>
<intersection>-28.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-28.5,40,-28.5</points>
<connection>
<GID>489</GID>
<name>IN_4</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-28,36.5,-28</points>
<connection>
<GID>491</GID>
<name>OUT_0</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>473 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-27.5,33,-26</points>
<intersection>-27.5 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-27.5,40,-27.5</points>
<connection>
<GID>489</GID>
<name>IN_5</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-26,33,-26</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>639 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,1,169,3.5</points>
<intersection>1 2</intersection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161.5,3.5,169,3.5</points>
<connection>
<GID>714</GID>
<name>IN_0</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>169,1,175.5,1</points>
<connection>
<GID>712</GID>
<name>IN_6</name></connection>
<intersection>169 0</intersection></hsegment></shape></wire>
<wire>
<ID>474 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-26.5,33.5,-24</points>
<intersection>-26.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-24,33.5,-24</points>
<connection>
<GID>524</GID>
<name>IN_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-26.5,40,-26.5</points>
<connection>
<GID>489</GID>
<name>IN_6</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>465 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-23.5,43,-20.5</points>
<connection>
<GID>489</GID>
<name>SEL_1</name></connection>
<connection>
<GID>501</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>631 </ID>
<shape>
<hsegment>
<ID>6</ID>
<points>176.5,7,177.5,7</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<intersection>177.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>177.5,4,177.5,7</points>
<connection>
<GID>712</GID>
<name>SEL_2</name></connection>
<intersection>7 6</intersection></vsegment></shape></wire>
<wire>
<ID>466 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-23.5,41,-20.5</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<intersection>-23.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>41,-23.5,42,-23.5</points>
<connection>
<GID>489</GID>
<name>SEL_2</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>705 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-46,-13.5,-43</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-13.5,-43,-13,-43</points>
<intersection>-13.5 0</intersection>
<intersection>-13 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-13,-43,-13,-40</points>
<connection>
<GID>742</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>497 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,13.5,74,14</points>
<intersection>13.5 1</intersection>
<intersection>14 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,13.5,75.5,13.5</points>
<connection>
<GID>559</GID>
<name>IN_1</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>73,14,74,14</points>
<connection>
<GID>585</GID>
<name>IN_0</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>704 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-46,-14.5,-43</points>
<connection>
<GID>490</GID>
<name>IN_1</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-15,-43,-14.5,-43</points>
<intersection>-15 3</intersection>
<intersection>-14.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-15,-43,-15,-40</points>
<connection>
<GID>759</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>703 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-46,-15.5,-43</points>
<connection>
<GID>490</GID>
<name>IN_2</name></connection>
<intersection>-43 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-16,-43,-16,-40</points>
<intersection>-43 2</intersection>
<intersection>-40 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-16,-43,-15.5,-43</points>
<intersection>-16 1</intersection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-17,-40,-16,-40</points>
<connection>
<GID>760</GID>
<name>IN_0</name></connection>
<intersection>-16 1</intersection></hsegment></shape></wire>
<wire>
<ID>702 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-46,-16.5,-43</points>
<connection>
<GID>490</GID>
<name>IN_3</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-19,-43,-16.5,-43</points>
<intersection>-19 3</intersection>
<intersection>-16.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-19,-43,-19,-40</points>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>709 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,-44.5,-3.5,-40</points>
<connection>
<GID>743</GID>
<name>IN_0</name></connection>
<intersection>-44.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-6.5,-46,-6.5,-44.5</points>
<connection>
<GID>490</GID>
<name>IN_B_0</name></connection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-6.5,-44.5,-3.5,-44.5</points>
<intersection>-6.5 1</intersection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>501 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,22,124.5,22.5</points>
<intersection>22 2</intersection>
<intersection>22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,22.5,131.5,22.5</points>
<connection>
<GID>637</GID>
<name>IN_3</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>117.5,22,124.5,22</points>
<connection>
<GID>791</GID>
<name>IN_0</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>708 </ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-7,-46,-7,-43</points>
<intersection>-46 3</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-7,-43,-5.5,-43</points>
<intersection>-7 1</intersection>
<intersection>-5.5 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-7.5,-46,-7,-46</points>
<connection>
<GID>490</GID>
<name>IN_B_1</name></connection>
<intersection>-7 1</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-5.5,-43,-5.5,-40</points>
<connection>
<GID>744</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>707 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8.5,-46,-8.5,-43</points>
<connection>
<GID>490</GID>
<name>IN_B_2</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-8.5,-43,-7.5,-43</points>
<intersection>-8.5 0</intersection>
<intersection>-7.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-7.5,-43,-7.5,-40</points>
<connection>
<GID>745</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>706 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-46,-9.5,-40</points>
<connection>
<GID>490</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>746</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>710 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-49.5,-2,-49</points>
<connection>
<GID>638</GID>
<name>OUT_0</name></connection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3.5,-49,-2,-49</points>
<connection>
<GID>490</GID>
<name>carry_in</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>725 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-55,-11,-54</points>
<connection>
<GID>490</GID>
<name>OUT_1</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-10.5,-56,-10.5,-55</points>
<connection>
<GID>644</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-11,-55,-10.5,-55</points>
<intersection>-11 0</intersection>
<intersection>-10.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>724 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-55,-12,-54</points>
<connection>
<GID>490</GID>
<name>OUT_2</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-12.5,-56,-12.5,-55</points>
<connection>
<GID>768</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-12.5,-55,-12,-55</points>
<intersection>-12.5 1</intersection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>649 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-34.5,170,-32</points>
<intersection>-34.5 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170,-32,175.5,-32</points>
<connection>
<GID>707</GID>
<name>IN_1</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161.5,-34.5,170,-34.5</points>
<connection>
<GID>730</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>472 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-28,29.5,-28</points>
<connection>
<GID>497</GID>
<name>IN_0</name></connection>
<connection>
<GID>491</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>573 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-8.5,119,-8</points>
<intersection>-8.5 2</intersection>
<intersection>-8 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>119,-8.5,120.5,-8.5</points>
<connection>
<GID>669</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>118,-8,119,-8</points>
<connection>
<GID>673</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>572 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-10.5,119,-10</points>
<intersection>-10.5 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-10.5,120.5,-10.5</points>
<connection>
<GID>669</GID>
<name>IN_1</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>118,-10,119,-10</points>
<connection>
<GID>640</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>402 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48,12.5,-48,12.5</points>
<connection>
<GID>804</GID>
<name>IN_4</name></connection>
<connection>
<GID>803</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>567 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-9.5,131.5,-4.5</points>
<intersection>-9.5 2</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,-4.5,132,-4.5</points>
<connection>
<GID>630</GID>
<name>IN_0</name></connection>
<intersection>131.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>126.5,-9.5,131.5,-9.5</points>
<connection>
<GID>669</GID>
<name>OUT</name></connection>
<intersection>131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>442 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,24,29,24</points>
<connection>
<GID>508</GID>
<name>IN_0</name></connection>
<connection>
<GID>492</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>467 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-38.5,27,-38</points>
<intersection>-38.5 1</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-38.5,28.5,-38.5</points>
<connection>
<GID>522</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-38,27,-38</points>
<connection>
<GID>499</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>734 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,5,-29,8.5</points>
<intersection>5 1</intersection>
<intersection>8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29,5,-27,5</points>
<connection>
<GID>777</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,8.5,-29,8.5</points>
<connection>
<GID>817</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>733 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,7,-28.5,9.5</points>
<intersection>7 1</intersection>
<intersection>9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-28.5,7,-27,7</points>
<connection>
<GID>778</GID>
<name>IN_0</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,9.5,-28.5,9.5</points>
<connection>
<GID>817</GID>
<name>IN_1</name></connection>
<intersection>-28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>731 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-29.5,11,-27,11</points>
<connection>
<GID>776</GID>
<name>IN_0</name></connection>
<intersection>-29.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-29.5,11,-29.5,11.5</points>
<connection>
<GID>817</GID>
<name>IN_3</name></connection>
<intersection>11 1</intersection></vsegment></shape></wire>
<wire>
<ID>730 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-29.5,13,-27,13</points>
<connection>
<GID>780</GID>
<name>IN_0</name></connection>
<intersection>-29.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-29.5,12.5,-29.5,13</points>
<connection>
<GID>817</GID>
<name>IN_4</name></connection>
<intersection>13 1</intersection></vsegment></shape></wire>
<wire>
<ID>729 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,13.5,-28,15</points>
<intersection>13.5 1</intersection>
<intersection>15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,13.5,-28,13.5</points>
<connection>
<GID>817</GID>
<name>IN_5</name></connection>
<intersection>-28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28,15,-27,15</points>
<connection>
<GID>781</GID>
<name>IN_0</name></connection>
<intersection>-28 0</intersection></hsegment></shape></wire>
<wire>
<ID>728 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,14.5,-29,17</points>
<intersection>14.5 2</intersection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29,17,-27,17</points>
<connection>
<GID>782</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,14.5,-29,14.5</points>
<connection>
<GID>817</GID>
<name>IN_6</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>727 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,15.5,-29.5,19</points>
<connection>
<GID>817</GID>
<name>IN_7</name></connection>
<intersection>19 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,19,-27,19</points>
<connection>
<GID>783</GID>
<name>IN_0</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>651 652 653 654 655 656 657 658 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36,12,-33.5,12</points>
<connection>
<GID>816</GID>
<name>OUT</name></connection>
<connection>
<GID>817</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>480 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-50.5,44,-47.5</points>
<connection>
<GID>529</GID>
<name>SEL_1</name></connection>
<connection>
<GID>541</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>620 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,19.5,168,21</points>
<intersection>19.5 1</intersection>
<intersection>21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161,19.5,168,19.5</points>
<connection>
<GID>704</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>168,21,175,21</points>
<connection>
<GID>678</GID>
<name>IN_2</name></connection>
<intersection>168 0</intersection></hsegment></shape></wire>
<wire>
<ID>665 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,-56,173,-55.5</points>
<intersection>-56 1</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173,-56,176.5,-56</points>
<connection>
<GID>733</GID>
<name>IN_4</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>170,-55.5,173,-55.5</points>
<connection>
<GID>734</GID>
<name>OUT_0</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>488 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-54.5,34,-53</points>
<intersection>-54.5 1</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-54.5,41,-54.5</points>
<connection>
<GID>529</GID>
<name>IN_5</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-53,34,-53</points>
<connection>
<GID>535</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>602 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-65.5,120,-65</points>
<intersection>-65.5 1</intersection>
<intersection>-65 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-65.5,121.5,-65.5</points>
<connection>
<GID>695</GID>
<name>IN_1</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>119,-65,120,-65</points>
<connection>
<GID>708</GID>
<name>IN_0</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>527 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-38.5,74.5,-38</points>
<intersection>-38.5 1</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-38.5,76,-38.5</points>
<connection>
<GID>601</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-38,74.5,-38</points>
<connection>
<GID>577</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>490 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-52.5,37,-51.5</points>
<connection>
<GID>503</GID>
<name>OUT_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-52.5,41,-52.5</points>
<connection>
<GID>529</GID>
<name>IN_7</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>601 </ID>
<shape>
<hsegment>
<ID>6</ID>
<points>134,-47.5,135,-47.5</points>
<connection>
<GID>675</GID>
<name>IN_0</name></connection>
<intersection>135 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>135,-50.5,135,-47.5</points>
<connection>
<GID>694</GID>
<name>SEL_2</name></connection>
<intersection>-47.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>424 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24,-12.5,-24,-10.5</points>
<connection>
<GID>506</GID>
<name>OUT_0</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,-12.5,-23,-12.5</points>
<connection>
<GID>504</GID>
<name>ENABLE</name></connection>
<intersection>-24 0</intersection></hsegment></shape></wire>
<wire>
<ID>593 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-27.5,125,-26</points>
<intersection>-27.5 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-27.5,132,-27.5</points>
<connection>
<GID>643</GID>
<name>IN_5</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>118,-26,125,-26</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>416 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,-14.5,-26.5,-8.5</points>
<intersection>-14.5 1</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-26.5,-14.5,-23,-14.5</points>
<connection>
<GID>504</GID>
<name>IN_7</name></connection>
<intersection>-26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-38,-8.5,-26.5,-8.5</points>
<connection>
<GID>505</GID>
<name>OUT_0</name></connection>
<intersection>-26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>478 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-55.5,37.5,-55</points>
<intersection>-55.5 1</intersection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-55.5,41,-55.5</points>
<connection>
<GID>529</GID>
<name>IN_4</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-55,37.5,-55</points>
<connection>
<GID>531</GID>
<name>OUT_0</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>627 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175,-10,175,-5</points>
<intersection>-10 2</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,-5,175.5,-5</points>
<connection>
<GID>712</GID>
<name>IN_0</name></connection>
<intersection>175 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>170,-10,175,-10</points>
<connection>
<GID>726</GID>
<name>OUT</name></connection>
<intersection>175 0</intersection></hsegment></shape></wire>
<wire>
<ID>634 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-6.5,170,-4</points>
<intersection>-6.5 2</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170,-4,175.5,-4</points>
<connection>
<GID>712</GID>
<name>IN_1</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161.5,-6.5,170,-6.5</points>
<connection>
<GID>713</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>486 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-57,81.5,-56.5</points>
<intersection>-57 2</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,-56.5,88.5,-56.5</points>
<connection>
<GID>609</GID>
<name>IN_3</name></connection>
<intersection>81.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-57,81.5,-57</points>
<connection>
<GID>790</GID>
<name>IN_0</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>635 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-4.5,168.5,-3</points>
<intersection>-4.5 1</intersection>
<intersection>-3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161.5,-4.5,168.5,-4.5</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<intersection>168.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>168.5,-3,175.5,-3</points>
<connection>
<GID>712</GID>
<name>IN_2</name></connection>
<intersection>168.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>576 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-2.5,168.5,-2</points>
<intersection>-2.5 2</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,-2,175.5,-2</points>
<connection>
<GID>712</GID>
<name>IN_3</name></connection>
<intersection>168.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161.5,-2.5,168.5,-2.5</points>
<connection>
<GID>796</GID>
<name>IN_0</name></connection>
<intersection>168.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>628 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172,-1,172,-0.5</points>
<intersection>-1 1</intersection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172,-1,175.5,-1</points>
<connection>
<GID>712</GID>
<name>IN_4</name></connection>
<intersection>172 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>169,-0.5,172,-0.5</points>
<connection>
<GID>696</GID>
<name>OUT_0</name></connection>
<intersection>172 0</intersection></hsegment></shape></wire>
<wire>
<ID>638 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,0,168.5,1.5</points>
<intersection>0 1</intersection>
<intersection>1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,0,175.5,0</points>
<connection>
<GID>712</GID>
<name>IN_5</name></connection>
<intersection>168.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161.5,1.5,168.5,1.5</points>
<connection>
<GID>543</GID>
<name>IN_0</name></connection>
<intersection>168.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>433 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,22,80,22.5</points>
<intersection>22 2</intersection>
<intersection>22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,22.5,87,22.5</points>
<connection>
<GID>557</GID>
<name>IN_3</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73,22,80,22</points>
<connection>
<GID>787</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>640 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171.5,2,171.5,3</points>
<connection>
<GID>711</GID>
<name>OUT_0</name></connection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171.5,2,175.5,2</points>
<connection>
<GID>712</GID>
<name>IN_7</name></connection>
<intersection>171.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>629 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,4,179.5,5.5</points>
<connection>
<GID>712</GID>
<name>SEL_0</name></connection>
<intersection>5.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>180.5,5.5,180.5,7</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<intersection>5.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>179.5,5.5,180.5,5.5</points>
<intersection>179.5 0</intersection>
<intersection>180.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>630 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,4,178.5,7</points>
<connection>
<GID>712</GID>
<name>SEL_1</name></connection>
<connection>
<GID>728</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>688 </ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-59.5,-46,-59.5,-43</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-59.5,-43,-59,-43</points>
<intersection>-59.5 1</intersection>
<intersection>-59 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-59,-43,-59,-40</points>
<connection>
<GID>764</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>689 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60.5,-46,-60.5,-43</points>
<connection>
<GID>507</GID>
<name>IN_1</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-61,-43,-60.5,-43</points>
<intersection>-61 3</intersection>
<intersection>-60.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-61,-43,-61,-40</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>687 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-61.5,-46,-61.5,-43</points>
<connection>
<GID>507</GID>
<name>IN_2</name></connection>
<intersection>-43 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-62,-43,-62,-40</points>
<intersection>-43 2</intersection>
<intersection>-40 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-62,-43,-61.5,-43</points>
<intersection>-62 1</intersection>
<intersection>-61.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-63,-40,-62,-40</points>
<connection>
<GID>765</GID>
<name>IN_0</name></connection>
<intersection>-62 1</intersection></hsegment></shape></wire>
<wire>
<ID>693 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52.5,-46,-52.5,-45</points>
<connection>
<GID>507</GID>
<name>IN_B_0</name></connection>
<intersection>-45 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-49,-45,-49,-40</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-52.5,-45,-49,-45</points>
<intersection>-52.5 0</intersection>
<intersection>-49 1</intersection></hsegment></shape></wire>
<wire>
<ID>692 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51,-44,-51,-40</points>
<connection>
<GID>752</GID>
<name>IN_0</name></connection>
<intersection>-44 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-53.5,-46,-53.5,-44</points>
<connection>
<GID>507</GID>
<name>IN_B_1</name></connection>
<intersection>-44 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-53.5,-44,-51,-44</points>
<intersection>-53.5 1</intersection>
<intersection>-51 0</intersection></hsegment></shape></wire>
<wire>
<ID>691 </ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-54.5,-46,-54.5,-43</points>
<connection>
<GID>507</GID>
<name>IN_B_2</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-54.5,-43,-53,-43</points>
<intersection>-54.5 1</intersection>
<intersection>-53 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-53,-43,-53,-40</points>
<connection>
<GID>753</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>690 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55.5,-46,-55.5,-43</points>
<connection>
<GID>507</GID>
<name>IN_B_3</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-55.5,-43,-55,-43</points>
<intersection>-55.5 0</intersection>
<intersection>-55 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-55,-43,-55,-40</points>
<connection>
<GID>754</GID>
<name>IN_0</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>718 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54.5,-56.5,-54.5,-55</points>
<connection>
<GID>771</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-56,-55,-56,-54</points>
<connection>
<GID>507</GID>
<name>OUT_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-56,-55,-54.5,-55</points>
<intersection>-56 1</intersection>
<intersection>-54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>717 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56.5,-56.5,-56.5,-55</points>
<connection>
<GID>656</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-57,-55,-57,-54</points>
<connection>
<GID>507</GID>
<name>OUT_1</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-57,-55,-56.5,-55</points>
<intersection>-57 1</intersection>
<intersection>-56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>509 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,4.5,91.5,6</points>
<connection>
<GID>550</GID>
<name>SEL_0</name></connection>
<intersection>6 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>92.5,6,92.5,7.5</points>
<connection>
<GID>597</GID>
<name>IN_0</name></connection>
<intersection>6 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>91.5,6,92.5,6</points>
<intersection>91.5 0</intersection>
<intersection>92.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>716 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58,-55,-58,-54</points>
<connection>
<GID>507</GID>
<name>OUT_2</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-58.5,-56.5,-58.5,-55</points>
<connection>
<GID>772</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-58.5,-55,-58,-55</points>
<intersection>-58.5 1</intersection>
<intersection>-58 0</intersection></hsegment></shape></wire>
<wire>
<ID>715 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60.5,-56.5,-60.5,-55</points>
<connection>
<GID>647</GID>
<name>IN_0</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-59,-55,-59,-54</points>
<connection>
<GID>507</GID>
<name>OUT_3</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-60.5,-55,-59,-55</points>
<intersection>-60.5 0</intersection>
<intersection>-59 1</intersection></hsegment></shape></wire>
<wire>
<ID>399 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48,8.5,-48,8.5</points>
<connection>
<GID>685</GID>
<name>IN_0</name></connection>
<connection>
<GID>804</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>547 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-55,78,-55</points>
<connection>
<GID>616</GID>
<name>IN_0</name></connection>
<connection>
<GID>611</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>398 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48,10.5,-48,10.5</points>
<connection>
<GID>685</GID>
<name>IN_2</name></connection>
<connection>
<GID>804</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>750 751 752 753 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60,-6,-60,10</points>
<intersection>-6 1</intersection>
<intersection>10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69.5,-6,-60,-6</points>
<connection>
<GID>593</GID>
<name>OUT</name></connection>
<intersection>-60 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-60,10,-52,10</points>
<connection>
<GID>685</GID>
<name>OUT</name></connection>
<intersection>-60 0</intersection></hsegment></shape></wire>
<wire>
<ID>662 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171.5,-26,171.5,-25</points>
<connection>
<GID>716</GID>
<name>OUT_0</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171.5,-26,175.5,-26</points>
<connection>
<GID>707</GID>
<name>IN_7</name></connection>
<intersection>171.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>487 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-55,30.5,-55</points>
<connection>
<GID>536</GID>
<name>IN_0</name></connection>
<connection>
<GID>531</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>491 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-56,47,-56</points>
<connection>
<GID>528</GID>
<name>IN_0</name></connection>
<connection>
<GID>529</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>477 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-64.5,40.5,-59.5</points>
<intersection>-64.5 2</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-59.5,41,-59.5</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-64.5,40.5,-64.5</points>
<connection>
<GID>530</GID>
<name>OUT</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>661 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,-27,169,-24.5</points>
<intersection>-27 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161.5,-24.5,169,-24.5</points>
<connection>
<GID>570</GID>
<name>IN_0</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>169,-27,175.5,-27</points>
<connection>
<GID>707</GID>
<name>IN_6</name></connection>
<intersection>169 0</intersection></hsegment></shape></wire>
<wire>
<ID>484 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-61,35.5,-58.5</points>
<intersection>-61 2</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-58.5,41,-58.5</points>
<connection>
<GID>529</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-61,35.5,-61</points>
<connection>
<GID>532</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>485 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-59,34,-57.5</points>
<intersection>-59 1</intersection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-59,34,-59</points>
<connection>
<GID>533</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-57.5,41,-57.5</points>
<connection>
<GID>529</GID>
<name>IN_2</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>609 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-53.5,126.5,-51</points>
<intersection>-53.5 2</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-51,126.5,-51</points>
<connection>
<GID>701</GID>
<name>IN_0</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>126.5,-53.5,133,-53.5</points>
<connection>
<GID>694</GID>
<name>IN_6</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>432 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-57,34,-56.5</points>
<intersection>-57 2</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-56.5,41,-56.5</points>
<connection>
<GID>529</GID>
<name>IN_3</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-57,34,-57</points>
<connection>
<GID>786</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>489 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-53.5,34.5,-51</points>
<intersection>-53.5 2</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-51,34.5,-51</points>
<connection>
<GID>534</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-53.5,41,-53.5</points>
<connection>
<GID>529</GID>
<name>IN_6</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>479 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-50.5,45,-49</points>
<connection>
<GID>529</GID>
<name>SEL_0</name></connection>
<intersection>-49 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>46,-49,46,-47.5</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<intersection>-49 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45,-49,46,-49</points>
<intersection>45 0</intersection>
<intersection>46 1</intersection></hsegment></shape></wire>
<wire>
<ID>481 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-50.5,42,-47.5</points>
<connection>
<GID>542</GID>
<name>IN_0</name></connection>
<intersection>-50.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>42,-50.5,43,-50.5</points>
<connection>
<GID>529</GID>
<name>SEL_2</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>483 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-63.5,28,-63</points>
<intersection>-63.5 2</intersection>
<intersection>-63 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28,-63.5,29.5,-63.5</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27,-63,28,-63</points>
<connection>
<GID>537</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>519 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,1.5,81,4</points>
<intersection>1.5 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,4,81,4</points>
<connection>
<GID>556</GID>
<name>IN_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81,1.5,87.5,1.5</points>
<connection>
<GID>550</GID>
<name>IN_6</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>482 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-65.5,28,-65</points>
<intersection>-65.5 1</intersection>
<intersection>-65 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-65.5,29.5,-65.5</points>
<connection>
<GID>530</GID>
<name>IN_1</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27,-65,28,-65</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>543 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-63.5,75.5,-63</points>
<intersection>-63.5 2</intersection>
<intersection>-63 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>75.5,-63.5,77,-63.5</points>
<connection>
<GID>610</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>74.5,-63,75.5,-63</points>
<connection>
<GID>617</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>506 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,23,93,23</points>
<connection>
<GID>545</GID>
<name>IN_0</name></connection>
<connection>
<GID>557</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>618 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,15,162,15.5</points>
<intersection>15 2</intersection>
<intersection>15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161,15.5,162,15.5</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162,15,163.5,15</points>
<connection>
<GID>715</GID>
<name>IN_0</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>520 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,2.5,83.5,3.5</points>
<connection>
<GID>547</GID>
<name>OUT_0</name></connection>
<intersection>2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,2.5,87.5,2.5</points>
<connection>
<GID>550</GID>
<name>IN_7</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>521 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-1,93.5,-1</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<connection>
<GID>550</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>624 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,25,168.5,27.5</points>
<intersection>25 2</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161,27.5,168.5,27.5</points>
<connection>
<GID>549</GID>
<name>IN_0</name></connection>
<intersection>168.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>168.5,25,175,25</points>
<connection>
<GID>678</GID>
<name>IN_6</name></connection>
<intersection>168.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>507 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-9.5,87,-4.5</points>
<intersection>-9.5 2</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-4.5,87.5,-4.5</points>
<connection>
<GID>550</GID>
<name>IN_0</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-9.5,87,-9.5</points>
<connection>
<GID>590</GID>
<name>OUT</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>514 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-6,82,-3.5</points>
<intersection>-6 2</intersection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-3.5,87.5,-3.5</points>
<connection>
<GID>550</GID>
<name>IN_1</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-6,82,-6</points>
<connection>
<GID>553</GID>
<name>IN_0</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>494 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,28.5,91,30</points>
<connection>
<GID>557</GID>
<name>SEL_0</name></connection>
<intersection>30 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>92,30,92,31.5</points>
<connection>
<GID>586</GID>
<name>IN_0</name></connection>
<intersection>30 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>91,30,92,30</points>
<intersection>91 0</intersection>
<intersection>92 1</intersection></hsegment></shape></wire>
<wire>
<ID>515 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-4,80.5,-2.5</points>
<intersection>-4 1</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-4,80.5,-4</points>
<connection>
<GID>554</GID>
<name>IN_0</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80.5,-2.5,87.5,-2.5</points>
<connection>
<GID>550</GID>
<name>IN_2</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>456 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-2,80.5,-1.5</points>
<intersection>-2 2</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-1.5,87.5,-1.5</points>
<connection>
<GID>550</GID>
<name>IN_3</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-2,80.5,-2</points>
<connection>
<GID>788</GID>
<name>IN_0</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>518 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,0.5,80.5,2</points>
<intersection>0.5 1</intersection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,0.5,87.5,0.5</points>
<connection>
<GID>550</GID>
<name>IN_5</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,2,80.5,2</points>
<connection>
<GID>591</GID>
<name>IN_0</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>511 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,4.5,88.5,7.5</points>
<connection>
<GID>599</GID>
<name>IN_0</name></connection>
<intersection>4.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>88.5,4.5,89.5,4.5</points>
<connection>
<GID>550</GID>
<name>SEL_2</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>517 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,0,77,0</points>
<connection>
<GID>594</GID>
<name>IN_0</name></connection>
<connection>
<GID>551</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>616 </ID>
<shape>
<hsegment>
<ID>6</ID>
<points>176,31,177,31</points>
<connection>
<GID>552</GID>
<name>IN_0</name></connection>
<intersection>177 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>177,28,177,31</points>
<connection>
<GID>678</GID>
<name>SEL_2</name></connection>
<intersection>31 6</intersection></vsegment></shape></wire>
<wire>
<ID>647 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162.5,-39,162.5,-38.5</points>
<intersection>-39 1</intersection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,-39,164,-39</points>
<connection>
<GID>555</GID>
<name>IN_1</name></connection>
<intersection>162.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>161.5,-38.5,162.5,-38.5</points>
<connection>
<GID>721</GID>
<name>IN_0</name></connection>
<intersection>162.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>642 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175,-38,175,-33</points>
<intersection>-38 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,-33,175.5,-33</points>
<connection>
<GID>707</GID>
<name>IN_0</name></connection>
<intersection>175 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>170,-38,175,-38</points>
<connection>
<GID>555</GID>
<name>OUT</name></connection>
<intersection>175 0</intersection></hsegment></shape></wire>
<wire>
<ID>669 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-66,163.5,-65.5</points>
<intersection>-66 1</intersection>
<intersection>-65.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163.5,-66,165,-66</points>
<connection>
<GID>581</GID>
<name>IN_1</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>162.5,-65.5,163.5,-65.5</points>
<connection>
<GID>738</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>492 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,14.5,86.5,19.5</points>
<intersection>14.5 2</intersection>
<intersection>19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,19.5,87,19.5</points>
<connection>
<GID>557</GID>
<name>IN_0</name></connection>
<intersection>86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,14.5,86.5,14.5</points>
<connection>
<GID>559</GID>
<name>OUT</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>499 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,18,81.5,20.5</points>
<intersection>18 2</intersection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,20.5,87,20.5</points>
<connection>
<GID>557</GID>
<name>IN_1</name></connection>
<intersection>81.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73,18,81.5,18</points>
<connection>
<GID>569</GID>
<name>IN_0</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>677 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182.5,-56.5,182.5,-56.5</points>
<connection>
<GID>567</GID>
<name>IN_0</name></connection>
<connection>
<GID>733</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>500 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,20,80,21.5</points>
<intersection>20 1</intersection>
<intersection>21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,20,80,20</points>
<connection>
<GID>572</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80,21.5,87,21.5</points>
<connection>
<GID>557</GID>
<name>IN_2</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>493 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,23.5,83.5,24</points>
<intersection>23.5 1</intersection>
<intersection>24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,23.5,87,23.5</points>
<connection>
<GID>557</GID>
<name>IN_4</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80.5,24,83.5,24</points>
<connection>
<GID>566</GID>
<name>OUT_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>503 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,24.5,80,26</points>
<intersection>24.5 1</intersection>
<intersection>26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,24.5,87,24.5</points>
<connection>
<GID>557</GID>
<name>IN_5</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73,26,80,26</points>
<connection>
<GID>578</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>495 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,28.5,90,31.5</points>
<connection>
<GID>557</GID>
<name>SEL_1</name></connection>
<connection>
<GID>588</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>673 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162.5,-55.5,166,-55.5</points>
<connection>
<GID>737</GID>
<name>IN_0</name></connection>
<connection>
<GID>734</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>496 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,28.5,88,31.5</points>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<intersection>28.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>88,28.5,89,28.5</points>
<connection>
<GID>557</GID>
<name>SEL_2</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>637 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>161.5,-0.5,165,-0.5</points>
<connection>
<GID>558</GID>
<name>IN_0</name></connection>
<connection>
<GID>696</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>535 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-25.5,83.5,-24.5</points>
<connection>
<GID>562</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-25.5,87.5,-25.5</points>
<connection>
<GID>563</GID>
<name>IN_7</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>498 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,15.5,74,16</points>
<intersection>15.5 2</intersection>
<intersection>16 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>74,15.5,75.5,15.5</points>
<connection>
<GID>559</GID>
<name>IN_0</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>73,16,74,16</points>
<connection>
<GID>583</GID>
<name>IN_0</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>512 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-10.5,74.5,-10</points>
<intersection>-10.5 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-10.5,76,-10.5</points>
<connection>
<GID>590</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-10,74.5,-10</points>
<connection>
<GID>560</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>614 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,28,179,29.5</points>
<connection>
<GID>678</GID>
<name>SEL_0</name></connection>
<intersection>29.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>180,29.5,180,31</points>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<intersection>29.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>179,29.5,180,29.5</points>
<intersection>179 0</intersection>
<intersection>180 1</intersection></hsegment></shape></wire>
<wire>
<ID>522 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-37.5,87,-32.5</points>
<intersection>-37.5 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-32.5,87.5,-32.5</points>
<connection>
<GID>563</GID>
<name>IN_0</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-37.5,87,-37.5</points>
<connection>
<GID>601</GID>
<name>OUT</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>529 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-34,82,-31.5</points>
<intersection>-34 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-31.5,87.5,-31.5</points>
<connection>
<GID>563</GID>
<name>IN_1</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-34,82,-34</points>
<connection>
<GID>602</GID>
<name>IN_0</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>530 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-32,80.5,-30.5</points>
<intersection>-32 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-32,80.5,-32</points>
<connection>
<GID>568</GID>
<name>IN_0</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80.5,-30.5,87.5,-30.5</points>
<connection>
<GID>563</GID>
<name>IN_2</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>471 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-30,80.5,-29.5</points>
<intersection>-30 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-29.5,87.5,-29.5</points>
<connection>
<GID>563</GID>
<name>IN_3</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-30,80.5,-30</points>
<connection>
<GID>789</GID>
<name>IN_0</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>502 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,24,76.5,24</points>
<connection>
<GID>582</GID>
<name>IN_0</name></connection>
<connection>
<GID>566</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>523 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-28.5,84,-28</points>
<intersection>-28.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-28.5,87.5,-28.5</points>
<connection>
<GID>563</GID>
<name>IN_4</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81,-28,84,-28</points>
<connection>
<GID>565</GID>
<name>OUT_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>533 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-27.5,80.5,-26</points>
<intersection>-27.5 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-27.5,87.5,-27.5</points>
<connection>
<GID>563</GID>
<name>IN_5</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-26,80.5,-26</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>534 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-26.5,81,-24</points>
<intersection>-26.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-24,81,-24</points>
<connection>
<GID>603</GID>
<name>IN_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81,-26.5,87.5,-26.5</points>
<connection>
<GID>563</GID>
<name>IN_6</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>524 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-23.5,91.5,-22</points>
<connection>
<GID>563</GID>
<name>SEL_0</name></connection>
<intersection>-22 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>92.5,-22,92.5,-20.5</points>
<connection>
<GID>605</GID>
<name>IN_0</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-22,92.5,-22</points>
<intersection>91.5 0</intersection>
<intersection>92.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>525 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-23.5,90.5,-20.5</points>
<connection>
<GID>563</GID>
<name>SEL_1</name></connection>
<connection>
<GID>579</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>526 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-23.5,88.5,-20.5</points>
<connection>
<GID>606</GID>
<name>IN_0</name></connection>
<intersection>-23.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>88.5,-23.5,89.5,-23.5</points>
<connection>
<GID>563</GID>
<name>SEL_2</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>536 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-29,93.5,-29</points>
<connection>
<GID>563</GID>
<name>OUT</name></connection>
<connection>
<GID>600</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>532 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-28,77,-28</points>
<connection>
<GID>574</GID>
<name>IN_0</name></connection>
<connection>
<GID>565</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>646 </ID>
<shape>
<hsegment>
<ID>6</ID>
<points>176.5,-21,177.5,-21</points>
<connection>
<GID>576</GID>
<name>IN_0</name></connection>
<intersection>177.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>177.5,-24,177.5,-21</points>
<connection>
<GID>707</GID>
<name>SEL_2</name></connection>
<intersection>-21 6</intersection></vsegment></shape></wire>
<wire>
<ID>670 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-64,163.5,-63.5</points>
<intersection>-64 2</intersection>
<intersection>-63.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>163.5,-64,165,-64</points>
<connection>
<GID>581</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>162.5,-63.5,163.5,-63.5</points>
<connection>
<GID>592</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>664 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,-65,176,-60</points>
<intersection>-65 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176,-60,176.5,-60</points>
<connection>
<GID>733</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>171,-65,176,-65</points>
<connection>
<GID>581</GID>
<name>OUT</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>675 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-54,170,-51.5</points>
<intersection>-54 2</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,-51.5,170,-51.5</points>
<connection>
<GID>587</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>170,-54,176.5,-54</points>
<connection>
<GID>733</GID>
<name>IN_6</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>513 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-8.5,74.5,-8</points>
<intersection>-8.5 2</intersection>
<intersection>-8 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-8.5,76,-8.5</points>
<connection>
<GID>590</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>73.5,-8,74.5,-8</points>
<connection>
<GID>596</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>409 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,12.5,-40,12.5</points>
<connection>
<GID>804</GID>
<name>OUT_4</name></connection>
<connection>
<GID>816</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>744 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75,-9,-75,-7.5</points>
<intersection>-9 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76,-9,-75,-9</points>
<connection>
<GID>800</GID>
<name>OUT_0</name></connection>
<intersection>-75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-75,-7.5,-73.5,-7.5</points>
<connection>
<GID>593</GID>
<name>IN_0</name></connection>
<intersection>-75 0</intersection></hsegment></shape></wire>
<wire>
<ID>743 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76,-6.5,-73.5,-6.5</points>
<connection>
<GID>593</GID>
<name>IN_1</name></connection>
<intersection>-76 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-76,-7,-76,-6.5</points>
<connection>
<GID>800</GID>
<name>OUT_1</name></connection>
<intersection>-6.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>742 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76,-5.5,-73.5,-5.5</points>
<connection>
<GID>593</GID>
<name>IN_2</name></connection>
<intersection>-76 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-76,-5.5,-76,-5</points>
<connection>
<GID>800</GID>
<name>OUT_2</name></connection>
<intersection>-5.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>741 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75,-4.5,-75,-3</points>
<intersection>-4.5 2</intersection>
<intersection>-3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76,-3,-75,-3</points>
<connection>
<GID>800</GID>
<name>OUT_3</name></connection>
<intersection>-75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-75,-4.5,-73.5,-4.5</points>
<connection>
<GID>593</GID>
<name>IN_3</name></connection>
<intersection>-75 0</intersection></hsegment></shape></wire>
<wire>
<ID>671 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-61.5,171,-59</points>
<intersection>-61.5 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171,-59,176.5,-59</points>
<connection>
<GID>733</GID>
<name>IN_1</name></connection>
<intersection>171 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-61.5,171,-61.5</points>
<connection>
<GID>595</GID>
<name>IN_0</name></connection>
<intersection>171 0</intersection></hsegment></shape></wire>
<wire>
<ID>528 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-36.5,74.5,-36</points>
<intersection>-36.5 2</intersection>
<intersection>-36 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-36.5,76,-36.5</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>73.5,-36,74.5,-36</points>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>550 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-52.5,84.5,-51.5</points>
<connection>
<GID>607</GID>
<name>OUT_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,-52.5,88.5,-52.5</points>
<connection>
<GID>609</GID>
<name>IN_7</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>551 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,-56,94.5,-56</points>
<connection>
<GID>608</GID>
<name>IN_0</name></connection>
<connection>
<GID>609</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>537 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-64.5,88,-59.5</points>
<intersection>-64.5 2</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-59.5,88.5,-59.5</points>
<connection>
<GID>609</GID>
<name>IN_0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83,-64.5,88,-64.5</points>
<connection>
<GID>610</GID>
<name>OUT</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>544 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-61,83,-58.5</points>
<intersection>-61 2</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-58.5,88.5,-58.5</points>
<connection>
<GID>609</GID>
<name>IN_1</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-61,83,-61</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>545 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-59,81.5,-57.5</points>
<intersection>-59 1</intersection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-59,81.5,-59</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<intersection>81.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,-57.5,88.5,-57.5</points>
<connection>
<GID>609</GID>
<name>IN_2</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>538 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-55.5,85,-55</points>
<intersection>-55.5 1</intersection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-55.5,88.5,-55.5</points>
<connection>
<GID>609</GID>
<name>IN_4</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-55,85,-55</points>
<connection>
<GID>611</GID>
<name>OUT_0</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>548 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-54.5,81.5,-53</points>
<intersection>-54.5 1</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,-54.5,88.5,-54.5</points>
<connection>
<GID>609</GID>
<name>IN_5</name></connection>
<intersection>81.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-53,81.5,-53</points>
<connection>
<GID>615</GID>
<name>IN_0</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>549 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-53.5,82,-51</points>
<intersection>-53.5 2</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-51,82,-51</points>
<connection>
<GID>614</GID>
<name>IN_0</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-53.5,88.5,-53.5</points>
<connection>
<GID>609</GID>
<name>IN_6</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>540 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-50.5,91.5,-47.5</points>
<connection>
<GID>609</GID>
<name>SEL_1</name></connection>
<connection>
<GID>621</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>541 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-50.5,89.5,-47.5</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<intersection>-50.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>89.5,-50.5,90.5,-50.5</points>
<connection>
<GID>609</GID>
<name>SEL_2</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>542 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-65.5,75.5,-65</points>
<intersection>-65.5 1</intersection>
<intersection>-65 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-65.5,77,-65.5</points>
<connection>
<GID>610</GID>
<name>IN_1</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>74.5,-65,75.5,-65</points>
<connection>
<GID>618</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>565 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,26.5,127.5,27.5</points>
<connection>
<GID>624</GID>
<name>OUT_0</name></connection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127.5,26.5,131.5,26.5</points>
<connection>
<GID>637</GID>
<name>IN_7</name></connection>
<intersection>127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>566 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,23,137.5,23</points>
<connection>
<GID>625</GID>
<name>IN_0</name></connection>
<connection>
<GID>637</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>404 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48,14.5,-48,14.5</points>
<connection>
<GID>804</GID>
<name>IN_6</name></connection>
<connection>
<GID>803</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>581 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-1,138,-1</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<connection>
<GID>630</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>574 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-6,126.5,-3.5</points>
<intersection>-6 2</intersection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126.5,-3.5,132,-3.5</points>
<connection>
<GID>630</GID>
<name>IN_1</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>118,-6,126.5,-6</points>
<connection>
<GID>633</GID>
<name>IN_0</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>410 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,15.5,-40,15.5</points>
<connection>
<GID>804</GID>
<name>OUT_7</name></connection>
<connection>
<GID>816</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>575 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-4,125,-2.5</points>
<intersection>-4 1</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-4,125,-4</points>
<connection>
<GID>634</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-2.5,132,-2.5</points>
<connection>
<GID>630</GID>
<name>IN_2</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>516 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-2,125,-1.5</points>
<intersection>-2 2</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-1.5,132,-1.5</points>
<connection>
<GID>630</GID>
<name>IN_3</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>118,-2,125,-2</points>
<connection>
<GID>792</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>578 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,0.5,125,2</points>
<intersection>0.5 1</intersection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,0.5,132,0.5</points>
<connection>
<GID>630</GID>
<name>IN_5</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>118,2,125,2</points>
<connection>
<GID>670</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>579 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,1.5,125.5,4</points>
<intersection>1.5 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,4,125.5,4</points>
<connection>
<GID>636</GID>
<name>IN_0</name></connection>
<intersection>125.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125.5,1.5,132,1.5</points>
<connection>
<GID>630</GID>
<name>IN_6</name></connection>
<intersection>125.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>569 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,4.5,136,6</points>
<connection>
<GID>630</GID>
<name>SEL_0</name></connection>
<intersection>6 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>137,6,137,7.5</points>
<connection>
<GID>674</GID>
<name>IN_0</name></connection>
<intersection>6 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>136,6,137,6</points>
<intersection>136 0</intersection>
<intersection>137 1</intersection></hsegment></shape></wire>
<wire>
<ID>570 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,4.5,135,7.5</points>
<connection>
<GID>630</GID>
<name>SEL_1</name></connection>
<connection>
<GID>676</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>560 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,20,124.5,21.5</points>
<intersection>20 1</intersection>
<intersection>21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,20,124.5,20</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,21.5,131.5,21.5</points>
<connection>
<GID>637</GID>
<name>IN_2</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>553 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,23.5,128,24</points>
<intersection>23.5 1</intersection>
<intersection>24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,23.5,131.5,23.5</points>
<connection>
<GID>637</GID>
<name>IN_4</name></connection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,24,128,24</points>
<connection>
<GID>646</GID>
<name>OUT_0</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>564 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,25.5,125,28</points>
<intersection>25.5 2</intersection>
<intersection>28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,28,125,28</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,25.5,131.5,25.5</points>
<connection>
<GID>637</GID>
<name>IN_6</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>406 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,10.5,-40,10.5</points>
<connection>
<GID>804</GID>
<name>OUT_2</name></connection>
<connection>
<GID>816</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>555 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,28.5,134.5,31.5</points>
<connection>
<GID>637</GID>
<name>SEL_1</name></connection>
<connection>
<GID>666</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>556 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,28.5,132.5,31.5</points>
<connection>
<GID>667</GID>
<name>IN_0</name></connection>
<intersection>28.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,28.5,133.5,28.5</points>
<connection>
<GID>637</GID>
<name>SEL_2</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>595 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-25.5,128,-24.5</points>
<connection>
<GID>642</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,-25.5,132,-25.5</points>
<connection>
<GID>643</GID>
<name>IN_7</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>403 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48,13.5,-48,13.5</points>
<connection>
<GID>804</GID>
<name>IN_5</name></connection>
<connection>
<GID>803</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>735 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45,6.5,-45,6.5</points>
<connection>
<GID>804</GID>
<name>clock</name></connection>
<connection>
<GID>775</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>636 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,8.5,-40,8.5</points>
<connection>
<GID>804</GID>
<name>OUT_0</name></connection>
<connection>
<GID>816</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>411 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,9.5,-40,9.5</points>
<connection>
<GID>804</GID>
<name>OUT_1</name></connection>
<connection>
<GID>816</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>589 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-34,126.5,-31.5</points>
<intersection>-34 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126.5,-31.5,132,-31.5</points>
<connection>
<GID>643</GID>
<name>IN_1</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>118,-34,126.5,-34</points>
<connection>
<GID>682</GID>
<name>IN_0</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>412 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,11.5,-40,11.5</points>
<connection>
<GID>804</GID>
<name>OUT_3</name></connection>
<connection>
<GID>816</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>407 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,14.5,-40,14.5</points>
<connection>
<GID>804</GID>
<name>OUT_6</name></connection>
<connection>
<GID>816</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>582 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-37.5,131.5,-32.5</points>
<intersection>-37.5 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,-32.5,132,-32.5</points>
<connection>
<GID>643</GID>
<name>IN_0</name></connection>
<intersection>131.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>126.5,-37.5,131.5,-37.5</points>
<connection>
<GID>680</GID>
<name>OUT</name></connection>
<intersection>131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>590 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-32,125,-30.5</points>
<intersection>-32 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-32,125,-32</points>
<connection>
<GID>648</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-30.5,132,-30.5</points>
<connection>
<GID>643</GID>
<name>IN_2</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>594 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-26.5,125.5,-24</points>
<intersection>-26.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-24,125.5,-24</points>
<connection>
<GID>683</GID>
<name>IN_0</name></connection>
<intersection>125.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125.5,-26.5,132,-26.5</points>
<connection>
<GID>643</GID>
<name>IN_6</name></connection>
<intersection>125.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>584 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-23.5,136,-22</points>
<connection>
<GID>643</GID>
<name>SEL_0</name></connection>
<intersection>-22 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>137,-22,137,-20.5</points>
<connection>
<GID>688</GID>
<name>IN_0</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>136,-22,137,-22</points>
<intersection>136 0</intersection>
<intersection>137 1</intersection></hsegment></shape></wire>
<wire>
<ID>586 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-23.5,133,-20.5</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<intersection>-23.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>133,-23.5,134,-23.5</points>
<connection>
<GID>643</GID>
<name>SEL_2</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>596 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-29,138,-29</points>
<connection>
<GID>643</GID>
<name>OUT</name></connection>
<connection>
<GID>679</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>626 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181,22.5,181,22.5</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<connection>
<GID>678</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>612 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174.5,14,174.5,19</points>
<intersection>14 2</intersection>
<intersection>19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174.5,19,175,19</points>
<connection>
<GID>678</GID>
<name>IN_0</name></connection>
<intersection>174.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>169.5,14,174.5,14</points>
<connection>
<GID>715</GID>
<name>OUT</name></connection>
<intersection>174.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>561 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,21.5,168,22</points>
<intersection>21.5 2</intersection>
<intersection>22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,22,175,22</points>
<connection>
<GID>678</GID>
<name>IN_3</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161,21.5,168,21.5</points>
<connection>
<GID>795</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment></shape></wire>
<wire>
<ID>625 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,26,171,27</points>
<connection>
<GID>710</GID>
<name>OUT_0</name></connection>
<intersection>26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171,26,175,26</points>
<connection>
<GID>678</GID>
<name>IN_7</name></connection>
<intersection>171 0</intersection></hsegment></shape></wire>
<wire>
<ID>588 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-36.5,119,-36</points>
<intersection>-36.5 2</intersection>
<intersection>-36 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>119,-36.5,120.5,-36.5</points>
<connection>
<GID>680</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>118,-36,119,-36</points>
<connection>
<GID>686</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>599 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-50.5,137,-49</points>
<connection>
<GID>694</GID>
<name>SEL_0</name></connection>
<intersection>-49 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>138,-49,138,-47.5</points>
<connection>
<GID>684</GID>
<name>IN_0</name></connection>
<intersection>-49 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>137,-49,138,-49</points>
<intersection>137 0</intersection>
<intersection>138 1</intersection></hsegment></shape></wire>
<wire>
<ID>610 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-52.5,129,-51.5</points>
<connection>
<GID>691</GID>
<name>OUT_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129,-52.5,133,-52.5</points>
<connection>
<GID>694</GID>
<name>IN_7</name></connection>
<intersection>129 0</intersection></hsegment></shape></wire>
<wire>
<ID>632 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162.5,-11,162.5,-10.5</points>
<intersection>-11 1</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,-11,164,-11</points>
<connection>
<GID>726</GID>
<name>IN_1</name></connection>
<intersection>162.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161.5,-10.5,162.5,-10.5</points>
<connection>
<GID>693</GID>
<name>IN_0</name></connection>
<intersection>162.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>604 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-61,127.5,-58.5</points>
<intersection>-61 2</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127.5,-58.5,133,-58.5</points>
<connection>
<GID>694</GID>
<name>IN_1</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119,-61,127.5,-61</points>
<connection>
<GID>698</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>598 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-55.5,129.5,-55</points>
<intersection>-55.5 1</intersection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-55.5,133,-55.5</points>
<connection>
<GID>694</GID>
<name>IN_4</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>126.5,-55,129.5,-55</points>
<connection>
<GID>697</GID>
<name>OUT_0</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>608 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-54.5,126,-53</points>
<intersection>-54.5 1</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,-54.5,133,-54.5</points>
<connection>
<GID>694</GID>
<name>IN_5</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119,-53,126,-53</points>
<connection>
<GID>702</GID>
<name>IN_0</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>600 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-50.5,136,-47.5</points>
<connection>
<GID>694</GID>
<name>SEL_1</name></connection>
<connection>
<GID>709</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>607 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-55,122.5,-55</points>
<connection>
<GID>705</GID>
<name>IN_0</name></connection>
<connection>
<GID>697</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>622 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161,23.5,164.5,23.5</points>
<connection>
<GID>723</GID>
<name>IN_0</name></connection>
<connection>
<GID>699</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>650 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-32.5,168.5,-31</points>
<intersection>-32.5 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161.5,-32.5,168.5,-32.5</points>
<connection>
<GID>718</GID>
<name>IN_0</name></connection>
<intersection>168.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>168.5,-31,175.5,-31</points>
<connection>
<GID>707</GID>
<name>IN_2</name></connection>
<intersection>168.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>591 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-30.5,168.5,-30</points>
<intersection>-30.5 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,-30,175.5,-30</points>
<connection>
<GID>707</GID>
<name>IN_3</name></connection>
<intersection>168.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161.5,-30.5,168.5,-30.5</points>
<connection>
<GID>797</GID>
<name>IN_0</name></connection>
<intersection>168.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>643 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172,-29,172,-28.5</points>
<intersection>-29 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172,-29,175.5,-29</points>
<connection>
<GID>707</GID>
<name>IN_4</name></connection>
<intersection>172 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>169,-28.5,172,-28.5</points>
<connection>
<GID>717</GID>
<name>OUT_0</name></connection>
<intersection>172 0</intersection></hsegment></shape></wire>
<wire>
<ID>660 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-28,168.5,-26.5</points>
<intersection>-28 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,-28,175.5,-28</points>
<connection>
<GID>707</GID>
<name>IN_5</name></connection>
<intersection>168.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161.5,-26.5,168.5,-26.5</points>
<connection>
<GID>719</GID>
<name>IN_0</name></connection>
<intersection>168.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>663 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-29.5,181.5,-29.5</points>
<connection>
<GID>707</GID>
<name>OUT</name></connection>
<connection>
<GID>729</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>659 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,-28.5,165,-28.5</points>
<connection>
<GID>720</GID>
<name>IN_0</name></connection>
<connection>
<GID>717</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>633 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162.5,-9,162.5,-8.5</points>
<intersection>-9 2</intersection>
<intersection>-8.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-9,164,-9</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<intersection>162.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>161.5,-8.5,162.5,-8.5</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<intersection>162.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>676 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172.5,-53,172.5,-52</points>
<connection>
<GID>732</GID>
<name>OUT_0</name></connection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172.5,-53,176.5,-53</points>
<connection>
<GID>733</GID>
<name>IN_7</name></connection>
<intersection>172.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>672 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-59.5,169.5,-58</points>
<intersection>-59.5 1</intersection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,-59.5,169.5,-59.5</points>
<connection>
<GID>735</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>169.5,-58,176.5,-58</points>
<connection>
<GID>733</GID>
<name>IN_2</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>674 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-55,169.5,-53.5</points>
<intersection>-55 1</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-55,176.5,-55</points>
<connection>
<GID>733</GID>
<name>IN_5</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-53.5,169.5,-53.5</points>
<connection>
<GID>736</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>666 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180.5,-51,180.5,-49.5</points>
<connection>
<GID>733</GID>
<name>SEL_0</name></connection>
<intersection>-49.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>181.5,-49.5,181.5,-48</points>
<connection>
<GID>739</GID>
<name>IN_0</name></connection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>180.5,-49.5,181.5,-49.5</points>
<intersection>180.5 0</intersection>
<intersection>181.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>667 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-51,179.5,-48</points>
<connection>
<GID>733</GID>
<name>SEL_1</name></connection>
<connection>
<GID>740</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>668 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177.5,-51,177.5,-48</points>
<connection>
<GID>741</GID>
<name>IN_0</name></connection>
<intersection>-51 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>177.5,-51,178.5,-51</points>
<connection>
<GID>733</GID>
<name>SEL_2</name></connection>
<intersection>177.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0.527039,37.9959,331.804,-124.083</PageViewport>
<gate>
<ID>882</ID>
<type>DA_FROM</type>
<position>61,-108</position>
<input>
<ID>IN_0</ID>1144 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin0</lparam></gate>
<gate>
<ID>818</ID>
<type>AA_LABEL</type>
<position>24.5,-133</position>
<gparam>LABEL_TEXT Instruction Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>826</ID>
<type>AA_LABEL</type>
<position>26.5,-21.5</position>
<gparam>LABEL_TEXT Address Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>819</ID>
<type>AI_RAM_12x16</type>
<position>117,10</position>
<input>
<ID>ADDRESS_0</ID>759 </input>
<input>
<ID>ADDRESS_1</ID>757 </input>
<input>
<ID>ADDRESS_10</ID>761 </input>
<input>
<ID>ADDRESS_11</ID>767 </input>
<input>
<ID>ADDRESS_2</ID>758 </input>
<input>
<ID>ADDRESS_3</ID>760 </input>
<input>
<ID>ADDRESS_4</ID>764 </input>
<input>
<ID>ADDRESS_5</ID>768 </input>
<input>
<ID>ADDRESS_6</ID>766 </input>
<input>
<ID>ADDRESS_7</ID>762 </input>
<input>
<ID>ADDRESS_8</ID>765 </input>
<input>
<ID>ADDRESS_9</ID>763 </input>
<input>
<ID>DATA_IN_0</ID>812 </input>
<input>
<ID>DATA_IN_1</ID>817 </input>
<input>
<ID>DATA_IN_10</ID>821 </input>
<input>
<ID>DATA_IN_11</ID>807 </input>
<input>
<ID>DATA_IN_12</ID>808 </input>
<input>
<ID>DATA_IN_13</ID>811 </input>
<input>
<ID>DATA_IN_14</ID>816 </input>
<input>
<ID>DATA_IN_15</ID>809 </input>
<input>
<ID>DATA_IN_2</ID>819 </input>
<input>
<ID>DATA_IN_3</ID>813 </input>
<input>
<ID>DATA_IN_4</ID>814 </input>
<input>
<ID>DATA_IN_5</ID>806 </input>
<input>
<ID>DATA_IN_6</ID>820 </input>
<input>
<ID>DATA_IN_7</ID>810 </input>
<input>
<ID>DATA_IN_8</ID>815 </input>
<input>
<ID>DATA_IN_9</ID>818 </input>
<output>
<ID>DATA_OUT_0</ID>812 </output>
<output>
<ID>DATA_OUT_1</ID>817 </output>
<output>
<ID>DATA_OUT_10</ID>821 </output>
<output>
<ID>DATA_OUT_11</ID>807 </output>
<output>
<ID>DATA_OUT_12</ID>808 </output>
<output>
<ID>DATA_OUT_13</ID>811 </output>
<output>
<ID>DATA_OUT_14</ID>816 </output>
<output>
<ID>DATA_OUT_15</ID>809 </output>
<output>
<ID>DATA_OUT_2</ID>819 </output>
<output>
<ID>DATA_OUT_3</ID>813 </output>
<output>
<ID>DATA_OUT_4</ID>814 </output>
<output>
<ID>DATA_OUT_5</ID>806 </output>
<output>
<ID>DATA_OUT_6</ID>820 </output>
<output>
<ID>DATA_OUT_7</ID>810 </output>
<output>
<ID>DATA_OUT_8</ID>815 </output>
<output>
<ID>DATA_OUT_9</ID>818 </output>
<input>
<ID>ENABLE_0</ID>1167 </input>
<input>
<ID>write_clock</ID>1143 </input>
<input>
<ID>write_enable</ID>1166 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:0 16640</lparam>
<lparam>Address:1 16671</lparam>
<lparam>Address:32 61568</lparam>
<lparam>Address:33 63488</lparam>
<lparam>Address:34 12352</lparam>
<lparam>Address:35 28674</lparam>
<lparam>Address:36 28673</lparam>
<lparam>Address:37 28676</lparam>
<lparam>Address:38 61952</lparam>
<lparam>Address:39 28704</lparam>
<lparam>Address:40 61696</lparam>
<lparam>Address:41 62464</lparam>
<lparam>Address:42 61504</lparam>
<lparam>Address:43 61696</lparam>
<lparam>Address:44 28704</lparam>
<lparam>Address:45 28673</lparam>
<lparam>Address:64 106</lparam>
<lparam>Address:80 8530</lparam>
<lparam>Address:81 4432</lparam>
<lparam>Address:82 32866</lparam>
<lparam>Address:83 53408</lparam>
<lparam>Address:84 28736</lparam>
<lparam>Address:85 28704</lparam>
<lparam>Address:86 29696</lparam>
<lparam>Address:87 29184</lparam>
<lparam>Address:88 28680</lparam>
<lparam>Address:89 28673</lparam>
<lparam>Address:90 28688</lparam>
<lparam>Address:91 28928</lparam>
<lparam>Address:92 62464</lparam>
<lparam>Address:93 28673</lparam>
<lparam>Address:94 28704</lparam>
<lparam>Address:95 62464</lparam>
<lparam>Address:96 28673</lparam>
<lparam>Address:98 269</lparam>
<lparam>Address:160 176</lparam>
<lparam>Address:176 84</lparam>
<lparam>Address:177 28928</lparam>
<lparam>Address:178 28800</lparam>
<lparam>Address:179 49328</lparam>
<lparam>Address:180 62464</lparam>
<lparam>Address:256 8528</lparam>
<lparam>Address:257 37201</lparam>
<lparam>Address:258 33106</lparam>
<lparam>Address:259 12800</lparam>
<lparam>Address:260 28673</lparam>
<lparam>Address:261 20787</lparam>
<lparam>Address:262 170</lparam>
<lparam>Address:263 30720</lparam>
<lparam>Address:264 29184</lparam>
<lparam>Address:265 28674</lparam>
<lparam>Address:266 28704</lparam>
<lparam>Address:267 28674</lparam>
<lparam>Address:268 28673</lparam>
<lparam>Address:269 28704</lparam>
<lparam>Address:270 28688</lparam>
<lparam>Address:271 28673</lparam>
<lparam>Address:272 30720</lparam>
<lparam>Address:273 29184</lparam>
<lparam>Address:274 28680</lparam>
<lparam>Address:275 28673</lparam>
<lparam>Address:276 12803</lparam>
<lparam>Address:277 61952</lparam>
<lparam>Address:278 16661</lparam>
<lparam>Address:279 63488</lparam>
<lparam>Address:280 62464</lparam>
<lparam>Address:281 12804</lparam>
<lparam>Address:282 61696</lparam>
<lparam>Address:283 16666</lparam>
<lparam>Address:284 8528</lparam>
<lparam>Address:285 62464</lparam>
<lparam>Address:286 16670</lparam>
<lparam>Address:287 12593</lparam>
<lparam>Address:288 28800</lparam>
<lparam>Address:289 12594</lparam>
<lparam>Address:290 61952</lparam>
<lparam>Address:291 16679</lparam>
<lparam>Address:292 63488</lparam>
<lparam>Address:293 62464</lparam>
<lparam>Address:294 12805</lparam>
<lparam>Address:295 61696</lparam>
<lparam>Address:296 16683</lparam>
<lparam>Address:297 8529</lparam>
<lparam>Address:298 62464</lparam>
<lparam>Address:299 8498</lparam>
<lparam>Address:300 28736</lparam>
<lparam>Address:301 8497</lparam>
<lparam>Address:302 61568</lparam>
<lparam>Address:303 49152</lparam>
<lparam>Address:304 28673</lparam>
<lparam>Address:308 41267</lparam>
<lparam>Address:309 29696</lparam>
<lparam>Address:310 28928</lparam>
<lparam>Address:311 28800</lparam>
<lparam>Address:312 12801</lparam>
<lparam>Address:313 28736</lparam>
<lparam>Address:314 28704</lparam>
<lparam>Address:315 12802</lparam>
<lparam>Address:316 24883</lparam>
<lparam>Address:317 49459</lparam>
<lparam>Address:336 25</lparam>
<lparam>Address:337 25</lparam>
<lparam>Address:338 25</lparam></gate>
<gate>
<ID>820</ID>
<type>AI_REGISTER12</type>
<position>68.5,-48.5</position>
<input>
<ID>IN_0</ID>996 </input>
<input>
<ID>IN_1</ID>992 </input>
<input>
<ID>IN_10</ID>991 </input>
<input>
<ID>IN_11</ID>1001 </input>
<input>
<ID>IN_2</ID>997 </input>
<input>
<ID>IN_3</ID>995 </input>
<input>
<ID>IN_4</ID>993 </input>
<input>
<ID>IN_5</ID>998 </input>
<input>
<ID>IN_6</ID>990 </input>
<input>
<ID>IN_7</ID>999 </input>
<input>
<ID>IN_8</ID>994 </input>
<input>
<ID>IN_9</ID>1000 </input>
<output>
<ID>OUT_0</ID>833 </output>
<output>
<ID>OUT_1</ID>834 </output>
<output>
<ID>OUT_10</ID>827 </output>
<output>
<ID>OUT_11</ID>830 </output>
<output>
<ID>OUT_2</ID>831 </output>
<output>
<ID>OUT_3</ID>832 </output>
<output>
<ID>OUT_4</ID>824 </output>
<output>
<ID>OUT_5</ID>823 </output>
<output>
<ID>OUT_6</ID>825 </output>
<output>
<ID>OUT_7</ID>826 </output>
<output>
<ID>OUT_8</ID>829 </output>
<output>
<ID>OUT_9</ID>828 </output>
<input>
<ID>clear</ID>1161 </input>
<input>
<ID>clock</ID>1143 </input>
<input>
<ID>count_enable</ID>1172 </input>
<input>
<ID>count_up</ID>1173 </input>
<input>
<ID>load</ID>1171 </input>
<gparam>VALUE_BOX -2.4,-0.8,2.4,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 261</lparam>
<lparam>INPUT_BITS 12</lparam>
<lparam>MAX_COUNT 4095</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>821</ID>
<type>AM_REGISTER16</type>
<position>68,-71.5</position>
<input>
<ID>IN_0</ID>1015 </input>
<input>
<ID>IN_1</ID>1024 </input>
<input>
<ID>IN_10</ID>1026 </input>
<input>
<ID>IN_11</ID>1020 </input>
<input>
<ID>IN_12</ID>1017 </input>
<input>
<ID>IN_13</ID>1018 </input>
<input>
<ID>IN_14</ID>1019 </input>
<input>
<ID>IN_15</ID>1028 </input>
<input>
<ID>IN_2</ID>1023 </input>
<input>
<ID>IN_3</ID>1022 </input>
<input>
<ID>IN_4</ID>1027 </input>
<input>
<ID>IN_5</ID>1014 </input>
<input>
<ID>IN_6</ID>1021 </input>
<input>
<ID>IN_7</ID>1013 </input>
<input>
<ID>IN_8</ID>1016 </input>
<input>
<ID>IN_9</ID>1025 </input>
<output>
<ID>OUT_0</ID>867 </output>
<output>
<ID>OUT_1</ID>871 </output>
<output>
<ID>OUT_10</ID>864 </output>
<output>
<ID>OUT_11</ID>870 </output>
<output>
<ID>OUT_12</ID>859 </output>
<output>
<ID>OUT_13</ID>860 </output>
<output>
<ID>OUT_14</ID>873 </output>
<output>
<ID>OUT_15</ID>874 </output>
<output>
<ID>OUT_2</ID>865 </output>
<output>
<ID>OUT_3</ID>866 </output>
<output>
<ID>OUT_4</ID>868 </output>
<output>
<ID>OUT_5</ID>862 </output>
<output>
<ID>OUT_6</ID>869 </output>
<output>
<ID>OUT_7</ID>872 </output>
<output>
<ID>OUT_8</ID>863 </output>
<output>
<ID>OUT_9</ID>861 </output>
<input>
<ID>clear</ID>1162 </input>
<input>
<ID>clock</ID>1143 </input>
<input>
<ID>count_enable</ID>1175 </input>
<input>
<ID>count_up</ID>1174 </input>
<input>
<ID>load</ID>1176 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>822</ID>
<type>AA_LABEL</type>
<position>26.5,-46</position>
<gparam>LABEL_TEXT Program Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>823</ID>
<type>AA_LABEL</type>
<position>29,-70.5</position>
<gparam>LABEL_TEXT Data Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>824</ID>
<type>AI_REGISTER12</type>
<position>68,-24</position>
<input>
<ID>IN_0</ID>1002 </input>
<input>
<ID>IN_1</ID>1005 </input>
<input>
<ID>IN_10</ID>1012 </input>
<input>
<ID>IN_11</ID>1011 </input>
<input>
<ID>IN_2</ID>1008 </input>
<input>
<ID>IN_3</ID>1006 </input>
<input>
<ID>IN_4</ID>1009 </input>
<input>
<ID>IN_5</ID>1010 </input>
<input>
<ID>IN_6</ID>1007 </input>
<input>
<ID>IN_7</ID>1003 </input>
<input>
<ID>IN_8</ID>1004 </input>
<input>
<ID>IN_9</ID>1190 </input>
<output>
<ID>OUT_0</ID>777 </output>
<output>
<ID>OUT_1</ID>779 </output>
<output>
<ID>OUT_10</ID>775 </output>
<output>
<ID>OUT_11</ID>771 </output>
<output>
<ID>OUT_2</ID>778 </output>
<output>
<ID>OUT_3</ID>780 </output>
<output>
<ID>OUT_4</ID>773 </output>
<output>
<ID>OUT_5</ID>772 </output>
<output>
<ID>OUT_6</ID>776 </output>
<output>
<ID>OUT_7</ID>770 </output>
<output>
<ID>OUT_8</ID>769 </output>
<output>
<ID>OUT_9</ID>774 </output>
<input>
<ID>clear</ID>1160 </input>
<input>
<ID>clock</ID>1143 </input>
<input>
<ID>count_enable</ID>1169 </input>
<input>
<ID>count_up</ID>1170 </input>
<input>
<ID>load</ID>1168 </input>
<gparam>VALUE_BOX -2.4,-0.8,2.4,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 261</lparam>
<lparam>INPUT_BITS 12</lparam>
<lparam>MAX_COUNT 4095</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>825</ID>
<type>DA_FROM</type>
<position>111,-12</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>827</ID>
<type>BX_16X1_BUS_END</type>
<position>113,-46.5</position>
<input>
<ID>Bus_in_0</ID>858 </input>
<input>
<ID>IN_1</ID>856 </input>
<input>
<ID>IN_10</ID>849 </input>
<input>
<ID>IN_11</ID>847 </input>
<input>
<ID>IN_2</ID>857 </input>
<input>
<ID>IN_3</ID>855 </input>
<input>
<ID>IN_4</ID>850 </input>
<input>
<ID>IN_5</ID>853 </input>
<input>
<ID>IN_6</ID>851 </input>
<input>
<ID>IN_7</ID>854 </input>
<input>
<ID>IN_8</ID>852 </input>
<input>
<ID>IN_9</ID>848 </input>
<input>
<ID>OUT</ID>1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>828</ID>
<type>AA_LABEL</type>
<position>110,24</position>
<gparam>LABEL_TEXT 4kx16 RAM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>829</ID>
<type>BX_16X1_BUS_END</type>
<position>112.5,-71.5</position>
<input>
<ID>Bus_in_0</ID>890 </input>
<input>
<ID>IN_1</ID>882 </input>
<input>
<ID>IN_10</ID>881 </input>
<input>
<ID>IN_11</ID>883 </input>
<input>
<ID>IN_12</ID>884 </input>
<input>
<ID>IN_13</ID>879 </input>
<input>
<ID>IN_14</ID>887 </input>
<input>
<ID>IN_15</ID>886 </input>
<input>
<ID>IN_2</ID>888 </input>
<input>
<ID>IN_3</ID>880 </input>
<input>
<ID>IN_4</ID>876 </input>
<input>
<ID>IN_5</ID>875 </input>
<input>
<ID>IN_6</ID>878 </input>
<input>
<ID>IN_7</ID>877 </input>
<input>
<ID>IN_8</ID>889 </input>
<input>
<ID>IN_9</ID>885 </input>
<input>
<ID>OUT</ID>1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>830</ID>
<type>DA_FROM</type>
<position>51,-107</position>
<input>
<ID>IN_0</ID>1145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin1</lparam></gate>
<gate>
<ID>831</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>106,-71.5</position>
<input>
<ID>ENABLE_0</ID>1188 </input>
<input>
<ID>IN_0</ID>867 </input>
<input>
<ID>IN_1</ID>871 </input>
<input>
<ID>IN_10</ID>864 </input>
<input>
<ID>IN_11</ID>870 </input>
<input>
<ID>IN_12</ID>859 </input>
<input>
<ID>IN_13</ID>860 </input>
<input>
<ID>IN_14</ID>873 </input>
<input>
<ID>IN_15</ID>874 </input>
<input>
<ID>IN_2</ID>865 </input>
<input>
<ID>IN_3</ID>866 </input>
<input>
<ID>IN_4</ID>868 </input>
<input>
<ID>IN_5</ID>862 </input>
<input>
<ID>IN_6</ID>869 </input>
<input>
<ID>IN_7</ID>872 </input>
<input>
<ID>IN_8</ID>863 </input>
<input>
<ID>IN_9</ID>861 </input>
<output>
<ID>OUT_0</ID>890 </output>
<output>
<ID>OUT_1</ID>882 </output>
<output>
<ID>OUT_10</ID>881 </output>
<output>
<ID>OUT_11</ID>883 </output>
<output>
<ID>OUT_12</ID>884 </output>
<output>
<ID>OUT_13</ID>879 </output>
<output>
<ID>OUT_14</ID>887 </output>
<output>
<ID>OUT_15</ID>886 </output>
<output>
<ID>OUT_2</ID>888 </output>
<output>
<ID>OUT_3</ID>880 </output>
<output>
<ID>OUT_4</ID>876 </output>
<output>
<ID>OUT_5</ID>875 </output>
<output>
<ID>OUT_6</ID>878 </output>
<output>
<ID>OUT_7</ID>877 </output>
<output>
<ID>OUT_8</ID>889 </output>
<output>
<ID>OUT_9</ID>885 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>832</ID>
<type>AA_LABEL</type>
<position>27.5,-99.5</position>
<gparam>LABEL_TEXT AC Accumulator</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>833</ID>
<type>DA_FROM</type>
<position>51,-105</position>
<input>
<ID>IN_0</ID>1159 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin3</lparam></gate>
<gate>
<ID>834</ID>
<type>BX_16X1_BUS_END</type>
<position>112.5,-100.5</position>
<input>
<ID>Bus_in_0</ID>922 </input>
<input>
<ID>IN_1</ID>914 </input>
<input>
<ID>IN_10</ID>913 </input>
<input>
<ID>IN_11</ID>915 </input>
<input>
<ID>IN_12</ID>916 </input>
<input>
<ID>IN_13</ID>911 </input>
<input>
<ID>IN_14</ID>919 </input>
<input>
<ID>IN_15</ID>918 </input>
<input>
<ID>IN_2</ID>920 </input>
<input>
<ID>IN_3</ID>912 </input>
<input>
<ID>IN_4</ID>908 </input>
<input>
<ID>IN_5</ID>907 </input>
<input>
<ID>IN_6</ID>910 </input>
<input>
<ID>IN_7</ID>909 </input>
<input>
<ID>IN_8</ID>921 </input>
<input>
<ID>IN_9</ID>917 </input>
<input>
<ID>OUT</ID>1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>835</ID>
<type>AA_LABEL</type>
<position>147.5,-193.5</position>
<gparam>LABEL_TEXT Output Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>836</ID>
<type>AM_REGISTER16</type>
<position>148.5,-178.5</position>
<input>
<ID>IN_0</ID>1067 </input>
<input>
<ID>IN_1</ID>1066 </input>
<input>
<ID>IN_10</ID>1063 </input>
<input>
<ID>IN_11</ID>1073 </input>
<input>
<ID>IN_12</ID>1075 </input>
<input>
<ID>IN_13</ID>1072 </input>
<input>
<ID>IN_14</ID>1076 </input>
<input>
<ID>IN_15</ID>1064 </input>
<input>
<ID>IN_2</ID>1074 </input>
<input>
<ID>IN_3</ID>1068 </input>
<input>
<ID>IN_4</ID>1061 </input>
<input>
<ID>IN_5</ID>1062 </input>
<input>
<ID>IN_6</ID>1069 </input>
<input>
<ID>IN_7</ID>1070 </input>
<input>
<ID>IN_8</ID>1071 </input>
<input>
<ID>IN_9</ID>1065 </input>
<output>
<ID>OUT_0</ID>1101 </output>
<output>
<ID>OUT_1</ID>1102 </output>
<output>
<ID>OUT_10</ID>1099 </output>
<output>
<ID>OUT_11</ID>1100 </output>
<output>
<ID>OUT_12</ID>1096 </output>
<output>
<ID>OUT_13</ID>1094 </output>
<output>
<ID>OUT_14</ID>1093 </output>
<output>
<ID>OUT_15</ID>1097 </output>
<output>
<ID>OUT_2</ID>1103 </output>
<output>
<ID>OUT_3</ID>1105 </output>
<output>
<ID>OUT_4</ID>1104 </output>
<output>
<ID>OUT_5</ID>1106 </output>
<output>
<ID>OUT_6</ID>1107 </output>
<output>
<ID>OUT_7</ID>1108 </output>
<output>
<ID>OUT_8</ID>1098 </output>
<output>
<ID>OUT_9</ID>1095 </output>
<input>
<ID>clear</ID>754 </input>
<input>
<ID>clock</ID>1143 </input>
<input>
<ID>count_enable</ID>1186 </input>
<input>
<ID>load</ID>1187 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>837</ID>
<type>BW_8X1_BUS_END</type>
<position>75,-22</position>
<input>
<ID>IN_0</ID>773 </input>
<input>
<ID>IN_1</ID>772 </input>
<input>
<ID>IN_2</ID>776 </input>
<input>
<ID>IN_3</ID>770 </input>
<input>
<ID>IN_4</ID>769 </input>
<input>
<ID>IN_5</ID>774 </input>
<input>
<ID>IN_6</ID>775 </input>
<input>
<ID>IN_7</ID>771 </input>
<input>
<ID>OUT</ID>781 782 783 784 785 786 787 788 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>838</ID>
<type>EE_VDD</type>
<position>40,15</position>
<output>
<ID>OUT_0</ID>988 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>839</ID>
<type>BV_4x1_BUS_END</type>
<position>75,-28</position>
<input>
<ID>IN_0</ID>777 </input>
<input>
<ID>IN_1</ID>779 </input>
<input>
<ID>IN_2</ID>778 </input>
<input>
<ID>IN_3</ID>780 </input>
<input>
<ID>OUT</ID>789 790 791 792 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>840</ID>
<type>CC_PULSE</type>
<position>32.5,4.5</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>841</ID>
<type>BV_4x1_BUS_END</type>
<position>88,6</position>
<input>
<ID>IN_0</ID>759 </input>
<input>
<ID>IN_1</ID>757 </input>
<input>
<ID>IN_2</ID>758 </input>
<input>
<ID>IN_3</ID>760 </input>
<input>
<ID>OUT</ID>789 790 791 792 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>842</ID>
<type>FF_GND</type>
<position>40,9</position>
<output>
<ID>OUT_0</ID>989 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>843</ID>
<type>BW_8X1_BUS_END</type>
<position>88,12</position>
<input>
<ID>IN_0</ID>764 </input>
<input>
<ID>IN_1</ID>768 </input>
<input>
<ID>IN_2</ID>766 </input>
<input>
<ID>IN_3</ID>762 </input>
<input>
<ID>IN_4</ID>765 </input>
<input>
<ID>IN_5</ID>763 </input>
<input>
<ID>IN_6</ID>761 </input>
<input>
<ID>IN_7</ID>767 </input>
<input>
<ID>OUT</ID>781 782 783 784 785 786 787 788 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>844</ID>
<type>DE_TO</type>
<position>46,10.5</position>
<input>
<ID>IN_0</ID>989 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>845</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>105.5,-22</position>
<input>
<ID>ENABLE_0</ID>801 </input>
<input>
<ID>IN_0</ID>796 </input>
<input>
<ID>IN_1</ID>795 </input>
<input>
<ID>IN_2</ID>799 </input>
<input>
<ID>IN_3</ID>793 </input>
<input>
<ID>IN_4</ID>798 </input>
<input>
<ID>IN_5</ID>797 </input>
<input>
<ID>IN_6</ID>794 </input>
<input>
<ID>IN_7</ID>800 </input>
<output>
<ID>OUT_0</ID>839 </output>
<output>
<ID>OUT_1</ID>840 </output>
<output>
<ID>OUT_2</ID>841 </output>
<output>
<ID>OUT_3</ID>842 </output>
<output>
<ID>OUT_4</ID>843 </output>
<output>
<ID>OUT_5</ID>844 </output>
<output>
<ID>OUT_6</ID>845 </output>
<output>
<ID>OUT_7</ID>846 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>846</ID>
<type>BX_16X1_BUS_END</type>
<position>56,-22</position>
<input>
<ID>Bus_in_0</ID>1002 </input>
<input>
<ID>IN_1</ID>1005 </input>
<input>
<ID>IN_10</ID>1012 </input>
<input>
<ID>IN_11</ID>1011 </input>
<input>
<ID>IN_2</ID>1008 </input>
<input>
<ID>IN_3</ID>1006 </input>
<input>
<ID>IN_4</ID>1009 </input>
<input>
<ID>IN_5</ID>1010 </input>
<input>
<ID>IN_6</ID>1007 </input>
<input>
<ID>IN_7</ID>1003 </input>
<input>
<ID>IN_8</ID>1004 </input>
<input>
<ID>IN_9</ID>1190 </input>
<input>
<ID>OUT</ID>1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>847</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>105.5,-29.5</position>
<input>
<ID>ENABLE_0</ID>801 </input>
<input>
<ID>IN_0</ID>802 </input>
<input>
<ID>IN_1</ID>805 </input>
<input>
<ID>IN_2</ID>803 </input>
<input>
<ID>IN_3</ID>804 </input>
<output>
<ID>OUT_0</ID>835 </output>
<output>
<ID>OUT_1</ID>836 </output>
<output>
<ID>OUT_2</ID>837 </output>
<output>
<ID>OUT_3</ID>838 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>848</ID>
<type>BX_16X1_BUS_END</type>
<position>56.5,-46.5</position>
<input>
<ID>Bus_in_0</ID>996 </input>
<input>
<ID>IN_1</ID>992 </input>
<input>
<ID>IN_10</ID>991 </input>
<input>
<ID>IN_11</ID>1001 </input>
<input>
<ID>IN_2</ID>997 </input>
<input>
<ID>IN_3</ID>995 </input>
<input>
<ID>IN_4</ID>993 </input>
<input>
<ID>IN_5</ID>998 </input>
<input>
<ID>IN_6</ID>990 </input>
<input>
<ID>IN_7</ID>999 </input>
<input>
<ID>IN_8</ID>994 </input>
<input>
<ID>IN_9</ID>1000 </input>
<input>
<ID>OUT</ID>1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>849</ID>
<type>BW_8X1_BUS_END</type>
<position>85.5,-22</position>
<input>
<ID>IN_0</ID>796 </input>
<input>
<ID>IN_1</ID>795 </input>
<input>
<ID>IN_2</ID>799 </input>
<input>
<ID>IN_3</ID>793 </input>
<input>
<ID>IN_4</ID>798 </input>
<input>
<ID>IN_5</ID>797 </input>
<input>
<ID>IN_6</ID>794 </input>
<input>
<ID>IN_7</ID>800 </input>
<input>
<ID>OUT</ID>781 782 783 784 785 786 787 788 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>850</ID>
<type>BX_16X1_BUS_END</type>
<position>56.5,-71.5</position>
<input>
<ID>Bus_in_0</ID>1015 </input>
<input>
<ID>IN_1</ID>1024 </input>
<input>
<ID>IN_10</ID>1026 </input>
<input>
<ID>IN_11</ID>1020 </input>
<input>
<ID>IN_12</ID>1017 </input>
<input>
<ID>IN_13</ID>1018 </input>
<input>
<ID>IN_14</ID>1019 </input>
<input>
<ID>IN_15</ID>1028 </input>
<input>
<ID>IN_2</ID>1023 </input>
<input>
<ID>IN_3</ID>1022 </input>
<input>
<ID>IN_4</ID>1027 </input>
<input>
<ID>IN_5</ID>1014 </input>
<input>
<ID>IN_6</ID>1021 </input>
<input>
<ID>IN_7</ID>1013 </input>
<input>
<ID>IN_8</ID>1016 </input>
<input>
<ID>IN_9</ID>1025 </input>
<input>
<ID>OUT</ID>1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>851</ID>
<type>BV_4x1_BUS_END</type>
<position>85.5,-29.5</position>
<input>
<ID>IN_0</ID>802 </input>
<input>
<ID>IN_1</ID>805 </input>
<input>
<ID>IN_2</ID>803 </input>
<input>
<ID>IN_3</ID>804 </input>
<input>
<ID>OUT</ID>789 790 791 792 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>852</ID>
<type>BX_16X1_BUS_END</type>
<position>117,-3</position>
<input>
<ID>Bus_in_0</ID>812 </input>
<input>
<ID>IN_1</ID>817 </input>
<input>
<ID>IN_10</ID>821 </input>
<input>
<ID>IN_11</ID>807 </input>
<input>
<ID>IN_12</ID>808 </input>
<input>
<ID>IN_13</ID>811 </input>
<input>
<ID>IN_14</ID>816 </input>
<input>
<ID>IN_15</ID>809 </input>
<input>
<ID>IN_2</ID>819 </input>
<input>
<ID>IN_3</ID>813 </input>
<input>
<ID>IN_4</ID>814 </input>
<input>
<ID>IN_5</ID>806 </input>
<input>
<ID>IN_6</ID>820 </input>
<input>
<ID>IN_7</ID>810 </input>
<input>
<ID>IN_8</ID>815 </input>
<input>
<ID>IN_9</ID>818 </input>
<input>
<ID>OUT</ID>1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>853</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>106,-52.5</position>
<input>
<ID>ENABLE_0</ID>822 </input>
<input>
<ID>IN_0</ID>833 </input>
<input>
<ID>IN_1</ID>834 </input>
<input>
<ID>IN_2</ID>831 </input>
<input>
<ID>IN_3</ID>832 </input>
<output>
<ID>OUT_0</ID>858 </output>
<output>
<ID>OUT_1</ID>856 </output>
<output>
<ID>OUT_2</ID>857 </output>
<output>
<ID>OUT_3</ID>855 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>854</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>106,-46.5</position>
<input>
<ID>ENABLE_0</ID>822 </input>
<input>
<ID>IN_0</ID>824 </input>
<input>
<ID>IN_1</ID>823 </input>
<input>
<ID>IN_2</ID>825 </input>
<input>
<ID>IN_3</ID>826 </input>
<input>
<ID>IN_4</ID>829 </input>
<input>
<ID>IN_5</ID>828 </input>
<input>
<ID>IN_6</ID>827 </input>
<input>
<ID>IN_7</ID>830 </input>
<output>
<ID>OUT_0</ID>850 </output>
<output>
<ID>OUT_1</ID>853 </output>
<output>
<ID>OUT_2</ID>851 </output>
<output>
<ID>OUT_3</ID>854 </output>
<output>
<ID>OUT_4</ID>852 </output>
<output>
<ID>OUT_5</ID>848 </output>
<output>
<ID>OUT_6</ID>849 </output>
<output>
<ID>OUT_7</ID>847 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>855</ID>
<type>BX_16X1_BUS_END</type>
<position>112.5,-23</position>
<input>
<ID>Bus_in_0</ID>835 </input>
<input>
<ID>IN_1</ID>836 </input>
<input>
<ID>IN_10</ID>845 </input>
<input>
<ID>IN_11</ID>846 </input>
<input>
<ID>IN_2</ID>837 </input>
<input>
<ID>IN_3</ID>838 </input>
<input>
<ID>IN_4</ID>839 </input>
<input>
<ID>IN_5</ID>840 </input>
<input>
<ID>IN_6</ID>841 </input>
<input>
<ID>IN_7</ID>842 </input>
<input>
<ID>IN_8</ID>843 </input>
<input>
<ID>IN_9</ID>844 </input>
<input>
<ID>OUT</ID>1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>856</ID>
<type>DA_FROM</type>
<position>61,-106</position>
<input>
<ID>IN_0</ID>1146 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin2</lparam></gate>
<gate>
<ID>857</ID>
<type>AM_REGISTER16</type>
<position>68,-100.5</position>
<input>
<ID>IN_0</ID>1144 </input>
<input>
<ID>IN_1</ID>1145 </input>
<input>
<ID>IN_10</ID>1150 </input>
<input>
<ID>IN_11</ID>1155 </input>
<input>
<ID>IN_12</ID>1151 </input>
<input>
<ID>IN_13</ID>1154 </input>
<input>
<ID>IN_14</ID>1152 </input>
<input>
<ID>IN_15</ID>1153 </input>
<input>
<ID>IN_2</ID>1146 </input>
<input>
<ID>IN_3</ID>1159 </input>
<input>
<ID>IN_4</ID>1147 </input>
<input>
<ID>IN_5</ID>1158 </input>
<input>
<ID>IN_6</ID>1148 </input>
<input>
<ID>IN_7</ID>1157 </input>
<input>
<ID>IN_8</ID>1149 </input>
<input>
<ID>IN_9</ID>1156 </input>
<output>
<ID>OUT_0</ID>899 </output>
<output>
<ID>OUT_1</ID>903 </output>
<output>
<ID>OUT_10</ID>896 </output>
<output>
<ID>OUT_11</ID>902 </output>
<output>
<ID>OUT_12</ID>891 </output>
<output>
<ID>OUT_13</ID>892 </output>
<output>
<ID>OUT_14</ID>905 </output>
<output>
<ID>OUT_15</ID>906 </output>
<output>
<ID>OUT_2</ID>897 </output>
<output>
<ID>OUT_3</ID>898 </output>
<output>
<ID>OUT_4</ID>900 </output>
<output>
<ID>OUT_5</ID>894 </output>
<output>
<ID>OUT_6</ID>901 </output>
<output>
<ID>OUT_7</ID>904 </output>
<output>
<ID>OUT_8</ID>895 </output>
<output>
<ID>OUT_9</ID>893 </output>
<input>
<ID>clear</ID>1163 </input>
<input>
<ID>clock</ID>1143 </input>
<input>
<ID>count_enable</ID>1178 </input>
<input>
<ID>count_up</ID>1179 </input>
<input>
<ID>load</ID>1177 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>858</ID>
<type>DA_FROM</type>
<position>61,-104</position>
<input>
<ID>IN_0</ID>1147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin4</lparam></gate>
<gate>
<ID>859</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>107,-100.5</position>
<input>
<ID>ENABLE_0</ID>755 </input>
<input>
<ID>IN_0</ID>899 </input>
<input>
<ID>IN_1</ID>903 </input>
<input>
<ID>IN_10</ID>896 </input>
<input>
<ID>IN_11</ID>902 </input>
<input>
<ID>IN_12</ID>891 </input>
<input>
<ID>IN_13</ID>892 </input>
<input>
<ID>IN_14</ID>905 </input>
<input>
<ID>IN_15</ID>906 </input>
<input>
<ID>IN_2</ID>897 </input>
<input>
<ID>IN_3</ID>898 </input>
<input>
<ID>IN_4</ID>900 </input>
<input>
<ID>IN_5</ID>894 </input>
<input>
<ID>IN_6</ID>901 </input>
<input>
<ID>IN_7</ID>904 </input>
<input>
<ID>IN_8</ID>895 </input>
<input>
<ID>IN_9</ID>893 </input>
<output>
<ID>OUT_0</ID>922 </output>
<output>
<ID>OUT_1</ID>914 </output>
<output>
<ID>OUT_10</ID>913 </output>
<output>
<ID>OUT_11</ID>915 </output>
<output>
<ID>OUT_12</ID>916 </output>
<output>
<ID>OUT_13</ID>911 </output>
<output>
<ID>OUT_14</ID>919 </output>
<output>
<ID>OUT_15</ID>918 </output>
<output>
<ID>OUT_2</ID>920 </output>
<output>
<ID>OUT_3</ID>912 </output>
<output>
<ID>OUT_4</ID>908 </output>
<output>
<ID>OUT_5</ID>907 </output>
<output>
<ID>OUT_6</ID>910 </output>
<output>
<ID>OUT_7</ID>909 </output>
<output>
<ID>OUT_8</ID>921 </output>
<output>
<ID>OUT_9</ID>917 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>860</ID>
<type>DA_FROM</type>
<position>51,-103</position>
<input>
<ID>IN_0</ID>1158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin5</lparam></gate>
<gate>
<ID>861</ID>
<type>AM_REGISTER16</type>
<position>68.5,-133.5</position>
<input>
<ID>IN_0</ID>1035 </input>
<input>
<ID>IN_1</ID>1029 </input>
<input>
<ID>IN_10</ID>1036 </input>
<input>
<ID>IN_11</ID>1043 </input>
<input>
<ID>IN_12</ID>1042 </input>
<input>
<ID>IN_13</ID>1041 </input>
<input>
<ID>IN_14</ID>1044 </input>
<input>
<ID>IN_15</ID>1040 </input>
<input>
<ID>IN_2</ID>1033 </input>
<input>
<ID>IN_3</ID>1037 </input>
<input>
<ID>IN_4</ID>1038 </input>
<input>
<ID>IN_5</ID>1039 </input>
<input>
<ID>IN_6</ID>1031 </input>
<input>
<ID>IN_7</ID>1030 </input>
<input>
<ID>IN_8</ID>1032 </input>
<input>
<ID>IN_9</ID>1034 </input>
<output>
<ID>OUT_0</ID>931 </output>
<output>
<ID>OUT_1</ID>935 </output>
<output>
<ID>OUT_10</ID>928 </output>
<output>
<ID>OUT_11</ID>934 </output>
<output>
<ID>OUT_12</ID>923 </output>
<output>
<ID>OUT_13</ID>924 </output>
<output>
<ID>OUT_14</ID>937 </output>
<output>
<ID>OUT_15</ID>938 </output>
<output>
<ID>OUT_2</ID>929 </output>
<output>
<ID>OUT_3</ID>930 </output>
<output>
<ID>OUT_4</ID>932 </output>
<output>
<ID>OUT_5</ID>926 </output>
<output>
<ID>OUT_6</ID>933 </output>
<output>
<ID>OUT_7</ID>936 </output>
<output>
<ID>OUT_8</ID>927 </output>
<output>
<ID>OUT_9</ID>925 </output>
<input>
<ID>clear</ID>1164 </input>
<input>
<ID>clock</ID>1143 </input>
<input>
<ID>count_enable</ID>1181 </input>
<input>
<ID>count_up</ID>1182 </input>
<input>
<ID>load</ID>1180 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 28673</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>862</ID>
<type>BX_16X1_BUS_END</type>
<position>113,-133.5</position>
<input>
<ID>Bus_in_0</ID>954 </input>
<input>
<ID>IN_1</ID>946 </input>
<input>
<ID>IN_10</ID>945 </input>
<input>
<ID>IN_11</ID>947 </input>
<input>
<ID>IN_12</ID>948 </input>
<input>
<ID>IN_13</ID>943 </input>
<input>
<ID>IN_14</ID>951 </input>
<input>
<ID>IN_15</ID>950 </input>
<input>
<ID>IN_2</ID>952 </input>
<input>
<ID>IN_3</ID>944 </input>
<input>
<ID>IN_4</ID>940 </input>
<input>
<ID>IN_5</ID>939 </input>
<input>
<ID>IN_6</ID>942 </input>
<input>
<ID>IN_7</ID>941 </input>
<input>
<ID>IN_8</ID>953 </input>
<input>
<ID>IN_9</ID>949 </input>
<input>
<ID>OUT</ID>1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>863</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>107.5,-133.5</position>
<input>
<ID>ENABLE_0</ID>756 </input>
<input>
<ID>IN_0</ID>931 </input>
<input>
<ID>IN_1</ID>935 </input>
<input>
<ID>IN_10</ID>928 </input>
<input>
<ID>IN_11</ID>934 </input>
<input>
<ID>IN_12</ID>923 </input>
<input>
<ID>IN_13</ID>924 </input>
<input>
<ID>IN_14</ID>937 </input>
<input>
<ID>IN_15</ID>938 </input>
<input>
<ID>IN_2</ID>929 </input>
<input>
<ID>IN_3</ID>930 </input>
<input>
<ID>IN_4</ID>932 </input>
<input>
<ID>IN_5</ID>926 </input>
<input>
<ID>IN_6</ID>933 </input>
<input>
<ID>IN_7</ID>936 </input>
<input>
<ID>IN_8</ID>927 </input>
<input>
<ID>IN_9</ID>925 </input>
<output>
<ID>OUT_0</ID>954 </output>
<output>
<ID>OUT_1</ID>946 </output>
<output>
<ID>OUT_10</ID>945 </output>
<output>
<ID>OUT_11</ID>947 </output>
<output>
<ID>OUT_12</ID>948 </output>
<output>
<ID>OUT_13</ID>943 </output>
<output>
<ID>OUT_14</ID>951 </output>
<output>
<ID>OUT_15</ID>950 </output>
<output>
<ID>OUT_2</ID>952 </output>
<output>
<ID>OUT_3</ID>944 </output>
<output>
<ID>OUT_4</ID>940 </output>
<output>
<ID>OUT_5</ID>939 </output>
<output>
<ID>OUT_6</ID>942 </output>
<output>
<ID>OUT_7</ID>941 </output>
<output>
<ID>OUT_8</ID>953 </output>
<output>
<ID>OUT_9</ID>949 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>864</ID>
<type>AM_REGISTER16</type>
<position>68.5,-160</position>
<input>
<ID>IN_0</ID>1045 </input>
<input>
<ID>IN_1</ID>1056 </input>
<input>
<ID>IN_10</ID>1048 </input>
<input>
<ID>IN_11</ID>1049 </input>
<input>
<ID>IN_12</ID>1055 </input>
<input>
<ID>IN_13</ID>1050 </input>
<input>
<ID>IN_14</ID>1059 </input>
<input>
<ID>IN_15</ID>1060 </input>
<input>
<ID>IN_2</ID>1047 </input>
<input>
<ID>IN_3</ID>1051 </input>
<input>
<ID>IN_4</ID>1046 </input>
<input>
<ID>IN_5</ID>1057 </input>
<input>
<ID>IN_6</ID>1052 </input>
<input>
<ID>IN_7</ID>1054 </input>
<input>
<ID>IN_8</ID>1053 </input>
<input>
<ID>IN_9</ID>1058 </input>
<output>
<ID>OUT_0</ID>963 </output>
<output>
<ID>OUT_1</ID>967 </output>
<output>
<ID>OUT_10</ID>960 </output>
<output>
<ID>OUT_11</ID>966 </output>
<output>
<ID>OUT_12</ID>955 </output>
<output>
<ID>OUT_13</ID>956 </output>
<output>
<ID>OUT_14</ID>969 </output>
<output>
<ID>OUT_15</ID>970 </output>
<output>
<ID>OUT_2</ID>961 </output>
<output>
<ID>OUT_3</ID>962 </output>
<output>
<ID>OUT_4</ID>964 </output>
<output>
<ID>OUT_5</ID>958 </output>
<output>
<ID>OUT_6</ID>965 </output>
<output>
<ID>OUT_7</ID>968 </output>
<output>
<ID>OUT_8</ID>959 </output>
<output>
<ID>OUT_9</ID>957 </output>
<input>
<ID>clear</ID>1165 </input>
<input>
<ID>clock</ID>1143 </input>
<input>
<ID>count_enable</ID>1184 </input>
<input>
<ID>count_up</ID>1185 </input>
<input>
<ID>load</ID>1183 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>865</ID>
<type>BX_16X1_BUS_END</type>
<position>113,-160</position>
<input>
<ID>Bus_in_0</ID>986 </input>
<input>
<ID>IN_1</ID>978 </input>
<input>
<ID>IN_10</ID>977 </input>
<input>
<ID>IN_11</ID>979 </input>
<input>
<ID>IN_12</ID>980 </input>
<input>
<ID>IN_13</ID>975 </input>
<input>
<ID>IN_14</ID>983 </input>
<input>
<ID>IN_15</ID>982 </input>
<input>
<ID>IN_2</ID>984 </input>
<input>
<ID>IN_3</ID>976 </input>
<input>
<ID>IN_4</ID>972 </input>
<input>
<ID>IN_5</ID>971 </input>
<input>
<ID>IN_6</ID>974 </input>
<input>
<ID>IN_7</ID>973 </input>
<input>
<ID>IN_8</ID>985 </input>
<input>
<ID>IN_9</ID>981 </input>
<input>
<ID>OUT</ID>1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>866</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>106,-160</position>
<input>
<ID>ENABLE_0</ID>1189 </input>
<input>
<ID>IN_0</ID>963 </input>
<input>
<ID>IN_1</ID>967 </input>
<input>
<ID>IN_10</ID>960 </input>
<input>
<ID>IN_11</ID>966 </input>
<input>
<ID>IN_12</ID>955 </input>
<input>
<ID>IN_13</ID>956 </input>
<input>
<ID>IN_14</ID>969 </input>
<input>
<ID>IN_15</ID>970 </input>
<input>
<ID>IN_2</ID>961 </input>
<input>
<ID>IN_3</ID>962 </input>
<input>
<ID>IN_4</ID>964 </input>
<input>
<ID>IN_5</ID>958 </input>
<input>
<ID>IN_6</ID>965 </input>
<input>
<ID>IN_7</ID>968 </input>
<input>
<ID>IN_8</ID>959 </input>
<input>
<ID>IN_9</ID>957 </input>
<output>
<ID>OUT_0</ID>986 </output>
<output>
<ID>OUT_1</ID>978 </output>
<output>
<ID>OUT_10</ID>977 </output>
<output>
<ID>OUT_11</ID>979 </output>
<output>
<ID>OUT_12</ID>980 </output>
<output>
<ID>OUT_13</ID>975 </output>
<output>
<ID>OUT_14</ID>983 </output>
<output>
<ID>OUT_15</ID>982 </output>
<output>
<ID>OUT_2</ID>984 </output>
<output>
<ID>OUT_3</ID>976 </output>
<output>
<ID>OUT_4</ID>972 </output>
<output>
<ID>OUT_5</ID>971 </output>
<output>
<ID>OUT_6</ID>974 </output>
<output>
<ID>OUT_7</ID>973 </output>
<output>
<ID>OUT_8</ID>985 </output>
<output>
<ID>OUT_9</ID>981 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>867</ID>
<type>AA_LABEL</type>
<position>25,-159</position>
<gparam>LABEL_TEXT Temporary Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>868</ID>
<type>DE_TO</type>
<position>47,4.5</position>
<input>
<ID>IN_0</ID>1192 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>869</ID>
<type>DE_TO</type>
<position>44,13.5</position>
<input>
<ID>IN_0</ID>988 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID vdd</lparam></gate>
<gate>
<ID>870</ID>
<type>BX_16X1_BUS_END</type>
<position>57.5,-133.5</position>
<input>
<ID>Bus_in_0</ID>1035 </input>
<input>
<ID>IN_1</ID>1029 </input>
<input>
<ID>IN_10</ID>1036 </input>
<input>
<ID>IN_11</ID>1043 </input>
<input>
<ID>IN_12</ID>1042 </input>
<input>
<ID>IN_13</ID>1041 </input>
<input>
<ID>IN_14</ID>1044 </input>
<input>
<ID>IN_15</ID>1040 </input>
<input>
<ID>IN_2</ID>1033 </input>
<input>
<ID>IN_3</ID>1037 </input>
<input>
<ID>IN_4</ID>1038 </input>
<input>
<ID>IN_5</ID>1039 </input>
<input>
<ID>IN_6</ID>1031 </input>
<input>
<ID>IN_7</ID>1030 </input>
<input>
<ID>IN_8</ID>1032 </input>
<input>
<ID>IN_9</ID>1034 </input>
<input>
<ID>OUT</ID>1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>871</ID>
<type>BX_16X1_BUS_END</type>
<position>57.5,-160</position>
<input>
<ID>Bus_in_0</ID>1045 </input>
<input>
<ID>IN_1</ID>1056 </input>
<input>
<ID>IN_10</ID>1048 </input>
<input>
<ID>IN_11</ID>1049 </input>
<input>
<ID>IN_12</ID>1055 </input>
<input>
<ID>IN_13</ID>1050 </input>
<input>
<ID>IN_14</ID>1059 </input>
<input>
<ID>IN_15</ID>1060 </input>
<input>
<ID>IN_2</ID>1047 </input>
<input>
<ID>IN_3</ID>1051 </input>
<input>
<ID>IN_4</ID>1046 </input>
<input>
<ID>IN_5</ID>1057 </input>
<input>
<ID>IN_6</ID>1052 </input>
<input>
<ID>IN_7</ID>1054 </input>
<input>
<ID>IN_8</ID>1053 </input>
<input>
<ID>IN_9</ID>1058 </input>
<input>
<ID>OUT</ID>1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>872</ID>
<type>BX_16X1_BUS_END</type>
<position>139.5,-178.5</position>
<input>
<ID>Bus_in_0</ID>1067 </input>
<input>
<ID>IN_1</ID>1066 </input>
<input>
<ID>IN_10</ID>1063 </input>
<input>
<ID>IN_11</ID>1073 </input>
<input>
<ID>IN_12</ID>1075 </input>
<input>
<ID>IN_13</ID>1072 </input>
<input>
<ID>IN_14</ID>1076 </input>
<input>
<ID>IN_15</ID>1064 </input>
<input>
<ID>IN_2</ID>1074 </input>
<input>
<ID>IN_3</ID>1068 </input>
<input>
<ID>IN_4</ID>1061 </input>
<input>
<ID>IN_5</ID>1062 </input>
<input>
<ID>IN_6</ID>1069 </input>
<input>
<ID>IN_7</ID>1070 </input>
<input>
<ID>IN_8</ID>1071 </input>
<input>
<ID>IN_9</ID>1065 </input>
<input>
<ID>OUT</ID>1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>873</ID>
<type>DA_FROM</type>
<position>102.5,-150</position>
<input>
<ID>IN_0</ID>1189 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID trBus</lparam></gate>
<gate>
<ID>874</ID>
<type>BW_8X1_BUS_END</type>
<position>156,-174.5</position>
<input>
<ID>IN_0</ID>1098 </input>
<input>
<ID>IN_1</ID>1095 </input>
<input>
<ID>IN_2</ID>1099 </input>
<input>
<ID>IN_3</ID>1100 </input>
<input>
<ID>IN_4</ID>1096 </input>
<input>
<ID>IN_5</ID>1094 </input>
<input>
<ID>IN_6</ID>1093 </input>
<input>
<ID>IN_7</ID>1097 </input>
<input>
<ID>OUT</ID>1109 1110 1111 1112 1113 1114 1115 1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>875</ID>
<type>BW_8X1_BUS_END</type>
<position>156,-182.5</position>
<input>
<ID>IN_0</ID>1101 </input>
<input>
<ID>IN_1</ID>1102 </input>
<input>
<ID>IN_2</ID>1103 </input>
<input>
<ID>IN_3</ID>1105 </input>
<input>
<ID>IN_4</ID>1104 </input>
<input>
<ID>IN_5</ID>1106 </input>
<input>
<ID>IN_6</ID>1107 </input>
<input>
<ID>IN_7</ID>1108 </input>
<input>
<ID>OUT</ID>1125 1126 1127 1128 1129 1130 1131 1132 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>876</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>169.5,-175</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1122 </input>
<input>
<ID>IN_2</ID>1117 </input>
<input>
<ID>IN_3</ID>1124 </input>
<input>
<ID>IN_4</ID>1121 </input>
<input>
<ID>IN_5</ID>1120 </input>
<input>
<ID>IN_6</ID>1118 </input>
<input>
<ID>IN_7</ID>1123 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>877</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>184,-175</position>
<input>
<ID>IN_0</ID>1133 </input>
<input>
<ID>IN_1</ID>1134 </input>
<input>
<ID>IN_2</ID>1135 </input>
<input>
<ID>IN_3</ID>1136 </input>
<input>
<ID>IN_4</ID>1137 </input>
<input>
<ID>IN_5</ID>1139 </input>
<input>
<ID>IN_6</ID>1138 </input>
<input>
<ID>IN_7</ID>1140 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>878</ID>
<type>BW_8X1_BUS_END</type>
<position>162.5,-174.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1122 </input>
<input>
<ID>IN_2</ID>1117 </input>
<input>
<ID>IN_3</ID>1124 </input>
<input>
<ID>IN_4</ID>1121 </input>
<input>
<ID>IN_5</ID>1120 </input>
<input>
<ID>IN_6</ID>1118 </input>
<input>
<ID>IN_7</ID>1123 </input>
<input>
<ID>OUT</ID>1109 1110 1111 1112 1113 1114 1115 1116 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>879</ID>
<type>BW_8X1_BUS_END</type>
<position>177,-174.5</position>
<input>
<ID>IN_0</ID>1133 </input>
<input>
<ID>IN_1</ID>1134 </input>
<input>
<ID>IN_2</ID>1135 </input>
<input>
<ID>IN_3</ID>1136 </input>
<input>
<ID>IN_4</ID>1137 </input>
<input>
<ID>IN_5</ID>1139 </input>
<input>
<ID>IN_6</ID>1138 </input>
<input>
<ID>IN_7</ID>1140 </input>
<input>
<ID>OUT</ID>1125 1126 1127 1128 1129 1130 1131 1132 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>880</ID>
<type>DA_FROM</type>
<position>113,-36</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>881</ID>
<type>DA_FROM</type>
<position>141.5,11.5</position>
<input>
<ID>IN_0</ID>1143 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>883</ID>
<type>DA_FROM</type>
<position>61,-102</position>
<input>
<ID>IN_0</ID>1148 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin6</lparam></gate>
<gate>
<ID>884</ID>
<type>DA_FROM</type>
<position>51,-101</position>
<input>
<ID>IN_0</ID>1157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin7</lparam></gate>
<gate>
<ID>885</ID>
<type>DA_FROM</type>
<position>61,-100</position>
<input>
<ID>IN_0</ID>1149 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin8</lparam></gate>
<gate>
<ID>886</ID>
<type>DA_FROM</type>
<position>51,-99</position>
<input>
<ID>IN_0</ID>1156 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin9</lparam></gate>
<gate>
<ID>887</ID>
<type>DA_FROM</type>
<position>61,-98</position>
<input>
<ID>IN_0</ID>1150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin10</lparam></gate>
<gate>
<ID>888</ID>
<type>DA_FROM</type>
<position>51,-97</position>
<input>
<ID>IN_0</ID>1155 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin11</lparam></gate>
<gate>
<ID>889</ID>
<type>DA_FROM</type>
<position>61,-96</position>
<input>
<ID>IN_0</ID>1151 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin12</lparam></gate>
<gate>
<ID>890</ID>
<type>DA_FROM</type>
<position>51,-95</position>
<input>
<ID>IN_0</ID>1154 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin13</lparam></gate>
<gate>
<ID>891</ID>
<type>DA_FROM</type>
<position>61,-94</position>
<input>
<ID>IN_0</ID>1152 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin14</lparam></gate>
<gate>
<ID>892</ID>
<type>DA_FROM</type>
<position>51,-93</position>
<input>
<ID>IN_0</ID>1153 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acin15</lparam></gate>
<gate>
<ID>893</ID>
<type>DA_FROM</type>
<position>64.5,-32.5</position>
<input>
<ID>IN_0</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrAR</lparam></gate>
<gate>
<ID>894</ID>
<type>DA_FROM</type>
<position>67.5,-57</position>
<input>
<ID>IN_0</ID>1161 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrPC</lparam></gate>
<gate>
<ID>895</ID>
<type>DA_FROM</type>
<position>66.5,-82.5</position>
<input>
<ID>IN_0</ID>1162 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrDR</lparam></gate>
<gate>
<ID>896</ID>
<type>DA_FROM</type>
<position>65,-112</position>
<input>
<ID>IN_0</ID>1163 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrAC</lparam></gate>
<gate>
<ID>897</ID>
<type>DA_FROM</type>
<position>66,-144</position>
<input>
<ID>IN_0</ID>1164 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrIR</lparam></gate>
<gate>
<ID>898</ID>
<type>DA_FROM</type>
<position>66.5,-173</position>
<input>
<ID>IN_0</ID>1165 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrTR</lparam></gate>
<gate>
<ID>899</ID>
<type>DA_FROM</type>
<position>141.5,9.5</position>
<input>
<ID>IN_0</ID>1166 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID write_memory</lparam></gate>
<gate>
<ID>900</ID>
<type>DA_FROM</type>
<position>141.5,7.5</position>
<input>
<ID>IN_0</ID>1167 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID read_memory</lparam></gate>
<gate>
<ID>901</ID>
<type>DE_TO</type>
<position>102.5,-13.5</position>
<input>
<ID>IN_0</ID>802 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ar0</lparam></gate>
<gate>
<ID>902</ID>
<type>DE_TO</type>
<position>101.5,-5.5</position>
<input>
<ID>IN_0</ID>805 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ar1</lparam></gate>
<gate>
<ID>903</ID>
<type>DE_TO</type>
<position>100.5,-13.5</position>
<input>
<ID>IN_0</ID>803 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ar2</lparam></gate>
<gate>
<ID>904</ID>
<type>DE_TO</type>
<position>99.5,-5.5</position>
<input>
<ID>IN_0</ID>804 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ar3</lparam></gate>
<gate>
<ID>905</ID>
<type>DE_TO</type>
<position>98.5,-13.5</position>
<input>
<ID>IN_0</ID>796 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ar4</lparam></gate>
<gate>
<ID>906</ID>
<type>DE_TO</type>
<position>97.5,-5.5</position>
<input>
<ID>IN_0</ID>795 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ar5</lparam></gate>
<gate>
<ID>907</ID>
<type>DE_TO</type>
<position>96.5,-13.5</position>
<input>
<ID>IN_0</ID>799 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ar6</lparam></gate>
<gate>
<ID>908</ID>
<type>DE_TO</type>
<position>95.5,-5.5</position>
<input>
<ID>IN_0</ID>793 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ar7</lparam></gate>
<gate>
<ID>909</ID>
<type>DE_TO</type>
<position>94.5,-13.5</position>
<input>
<ID>IN_0</ID>798 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ar8</lparam></gate>
<gate>
<ID>910</ID>
<type>DE_TO</type>
<position>93.5,-5.5</position>
<input>
<ID>IN_0</ID>797 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ar9</lparam></gate>
<gate>
<ID>911</ID>
<type>DE_TO</type>
<position>92.5,-13.5</position>
<input>
<ID>IN_0</ID>794 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ar10</lparam></gate>
<gate>
<ID>912</ID>
<type>DE_TO</type>
<position>91.5,-5.5</position>
<input>
<ID>IN_0</ID>800 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ar11</lparam></gate>
<gate>
<ID>913</ID>
<type>DE_TO</type>
<position>103.5,-61.5</position>
<input>
<ID>IN_0</ID>867 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr0</lparam></gate>
<gate>
<ID>914</ID>
<type>DE_TO</type>
<position>101.5,-61.5</position>
<input>
<ID>IN_0</ID>871 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr1</lparam></gate>
<gate>
<ID>915</ID>
<type>DE_TO</type>
<position>99.5,-61.5</position>
<input>
<ID>IN_0</ID>865 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr2</lparam></gate>
<gate>
<ID>916</ID>
<type>DE_TO</type>
<position>97.5,-61.5</position>
<input>
<ID>IN_0</ID>866 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr3</lparam></gate>
<gate>
<ID>917</ID>
<type>DE_TO</type>
<position>95.5,-61.5</position>
<input>
<ID>IN_0</ID>868 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr4</lparam></gate>
<gate>
<ID>918</ID>
<type>DE_TO</type>
<position>93.5,-61.5</position>
<input>
<ID>IN_0</ID>862 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr5</lparam></gate>
<gate>
<ID>919</ID>
<type>DE_TO</type>
<position>91.5,-61.5</position>
<input>
<ID>IN_0</ID>869 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr6</lparam></gate>
<gate>
<ID>920</ID>
<type>DE_TO</type>
<position>89.5,-61.5</position>
<input>
<ID>IN_0</ID>872 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr7</lparam></gate>
<gate>
<ID>921</ID>
<type>DE_TO</type>
<position>87.5,-61.5</position>
<input>
<ID>IN_0</ID>863 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr8</lparam></gate>
<gate>
<ID>922</ID>
<type>DE_TO</type>
<position>85.5,-61.5</position>
<input>
<ID>IN_0</ID>861 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr9</lparam></gate>
<gate>
<ID>923</ID>
<type>DE_TO</type>
<position>83.5,-61.5</position>
<input>
<ID>IN_0</ID>864 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr10</lparam></gate>
<gate>
<ID>924</ID>
<type>DE_TO</type>
<position>81.5,-61.5</position>
<input>
<ID>IN_0</ID>870 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr11</lparam></gate>
<gate>
<ID>925</ID>
<type>DE_TO</type>
<position>79.5,-61.5</position>
<input>
<ID>IN_0</ID>859 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr12</lparam></gate>
<gate>
<ID>926</ID>
<type>DE_TO</type>
<position>77.5,-61.5</position>
<input>
<ID>IN_0</ID>860 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr13</lparam></gate>
<gate>
<ID>927</ID>
<type>DE_TO</type>
<position>75.5,-61.5</position>
<input>
<ID>IN_0</ID>873 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr14</lparam></gate>
<gate>
<ID>928</ID>
<type>DE_TO</type>
<position>73.5,-61.5</position>
<input>
<ID>IN_0</ID>874 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID dr15</lparam></gate>
<gate>
<ID>929</ID>
<type>DE_TO</type>
<position>104,-89</position>
<input>
<ID>IN_0</ID>899 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>930</ID>
<type>DE_TO</type>
<position>102,-89</position>
<input>
<ID>IN_0</ID>903 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>931</ID>
<type>DE_TO</type>
<position>100,-89</position>
<input>
<ID>IN_0</ID>897 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>932</ID>
<type>DE_TO</type>
<position>98,-89</position>
<input>
<ID>IN_0</ID>898 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>933</ID>
<type>DE_TO</type>
<position>96,-89</position>
<input>
<ID>IN_0</ID>900 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>934</ID>
<type>DE_TO</type>
<position>94,-89</position>
<input>
<ID>IN_0</ID>894 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>935</ID>
<type>DE_TO</type>
<position>92,-89</position>
<input>
<ID>IN_0</ID>901 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>936</ID>
<type>DE_TO</type>
<position>90,-89</position>
<input>
<ID>IN_0</ID>904 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>937</ID>
<type>DE_TO</type>
<position>88,-89</position>
<input>
<ID>IN_0</ID>895 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>938</ID>
<type>DE_TO</type>
<position>86,-89</position>
<input>
<ID>IN_0</ID>893 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>939</ID>
<type>DE_TO</type>
<position>84,-89</position>
<input>
<ID>IN_0</ID>896 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>940</ID>
<type>DA_FROM</type>
<position>59.5,-58.5</position>
<input>
<ID>IN_0</ID>1174 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID vdd</lparam></gate>
<gate>
<ID>941</ID>
<type>DE_TO</type>
<position>82,-89</position>
<input>
<ID>IN_0</ID>902 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>942</ID>
<type>DE_TO</type>
<position>80,-89</position>
<input>
<ID>IN_0</ID>891 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>943</ID>
<type>DE_TO</type>
<position>78,-89</position>
<input>
<ID>IN_0</ID>892 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>944</ID>
<type>DE_TO</type>
<position>76,-89</position>
<input>
<ID>IN_0</ID>905 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>945</ID>
<type>DE_TO</type>
<position>74,-89</position>
<input>
<ID>IN_0</ID>906 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>946</ID>
<type>DA_FROM</type>
<position>59.5,-62.5</position>
<input>
<ID>IN_0</ID>1176 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldDR</lparam></gate>
<gate>
<ID>947</ID>
<type>DE_TO</type>
<position>104.5,-122.5</position>
<input>
<ID>IN_0</ID>931 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir0</lparam></gate>
<gate>
<ID>948</ID>
<type>DE_TO</type>
<position>102.5,-122.5</position>
<input>
<ID>IN_0</ID>935 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir1</lparam></gate>
<gate>
<ID>949</ID>
<type>DA_FROM</type>
<position>61.5,-148</position>
<input>
<ID>IN_0</ID>1184 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incTR</lparam></gate>
<gate>
<ID>950</ID>
<type>DE_TO</type>
<position>100.5,-122.5</position>
<input>
<ID>IN_0</ID>929 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir2</lparam></gate>
<gate>
<ID>951</ID>
<type>DE_TO</type>
<position>98.5,-122.5</position>
<input>
<ID>IN_0</ID>930 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir3</lparam></gate>
<gate>
<ID>952</ID>
<type>DA_FROM</type>
<position>61.5,-88.5</position>
<input>
<ID>IN_0</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incAC</lparam></gate>
<gate>
<ID>953</ID>
<type>DE_TO</type>
<position>96.5,-122.5</position>
<input>
<ID>IN_0</ID>932 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir4</lparam></gate>
<gate>
<ID>954</ID>
<type>DE_TO</type>
<position>94.5,-122.5</position>
<input>
<ID>IN_0</ID>926 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir5</lparam></gate>
<gate>
<ID>955</ID>
<type>DA_FROM</type>
<position>64.5,-38</position>
<input>
<ID>IN_0</ID>1172 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incPC</lparam></gate>
<gate>
<ID>956</ID>
<type>DE_TO</type>
<position>92.5,-122.5</position>
<input>
<ID>IN_0</ID>933 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir6</lparam></gate>
<gate>
<ID>957</ID>
<type>DE_TO</type>
<position>90.5,-122.5</position>
<input>
<ID>IN_0</ID>936 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir7</lparam></gate>
<gate>
<ID>958</ID>
<type>DA_FROM</type>
<position>63.5,-118.5</position>
<input>
<ID>IN_0</ID>1182 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID vdd</lparam></gate>
<gate>
<ID>959</ID>
<type>DE_TO</type>
<position>88.5,-122.5</position>
<input>
<ID>IN_0</ID>927 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir8</lparam></gate>
<gate>
<ID>960</ID>
<type>DE_TO</type>
<position>86.5,-122.5</position>
<input>
<ID>IN_0</ID>925 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir9</lparam></gate>
<gate>
<ID>961</ID>
<type>DA_FROM</type>
<position>103,-40.5</position>
<input>
<ID>IN_0</ID>822 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID pcBus</lparam></gate>
<gate>
<ID>962</ID>
<type>DE_TO</type>
<position>84.5,-122.5</position>
<input>
<ID>IN_0</ID>928 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir10</lparam></gate>
<gate>
<ID>963</ID>
<type>DE_TO</type>
<position>82.5,-122.5</position>
<input>
<ID>IN_0</ID>934 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir11</lparam></gate>
<gate>
<ID>964</ID>
<type>DE_TO</type>
<position>80.5,-122.5</position>
<input>
<ID>IN_0</ID>923 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir12</lparam></gate>
<gate>
<ID>965</ID>
<type>DE_TO</type>
<position>78.5,-122.5</position>
<input>
<ID>IN_0</ID>924 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir13</lparam></gate>
<gate>
<ID>966</ID>
<type>DA_FROM</type>
<position>63.5,-122.5</position>
<input>
<ID>IN_0</ID>1180 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldIR</lparam></gate>
<gate>
<ID>967</ID>
<type>DE_TO</type>
<position>76.5,-122.5</position>
<input>
<ID>IN_0</ID>937 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir14</lparam></gate>
<gate>
<ID>968</ID>
<type>DE_TO</type>
<position>74.5,-122.5</position>
<input>
<ID>IN_0</ID>938 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ir15</lparam></gate>
<gate>
<ID>969</ID>
<type>DA_FROM</type>
<position>64.5,-15.5</position>
<input>
<ID>IN_0</ID>1168 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldAR</lparam></gate>
<gate>
<ID>970</ID>
<type>DA_FROM</type>
<position>64.5,-13.5</position>
<input>
<ID>IN_0</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incAR</lparam></gate>
<gate>
<ID>971</ID>
<type>DA_FROM</type>
<position>64.5,-11.5</position>
<input>
<ID>IN_0</ID>1170 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID vdd</lparam></gate>
<gate>
<ID>972</ID>
<type>DA_FROM</type>
<position>64.5,-40</position>
<input>
<ID>IN_0</ID>1171 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldPC</lparam></gate>
<gate>
<ID>973</ID>
<type>DA_FROM</type>
<position>64.5,-35.5</position>
<input>
<ID>IN_0</ID>1173 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID vdd</lparam></gate>
<gate>
<ID>974</ID>
<type>DA_FROM</type>
<position>59.5,-60.5</position>
<input>
<ID>IN_0</ID>1175 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incDR</lparam></gate>
<gate>
<ID>975</ID>
<type>DA_FROM</type>
<position>61.5,-90.5</position>
<input>
<ID>IN_0</ID>1177 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldAC</lparam></gate>
<gate>
<ID>976</ID>
<type>DA_FROM</type>
<position>61.5,-86.5</position>
<input>
<ID>IN_0</ID>1179 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID vdd</lparam></gate>
<gate>
<ID>977</ID>
<type>DA_FROM</type>
<position>63.5,-120.5</position>
<input>
<ID>IN_0</ID>1181 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incIR</lparam></gate>
<gate>
<ID>978</ID>
<type>DA_FROM</type>
<position>61.5,-150</position>
<input>
<ID>IN_0</ID>1183 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldTR</lparam></gate>
<gate>
<ID>979</ID>
<type>DA_FROM</type>
<position>61.5,-146</position>
<input>
<ID>IN_0</ID>1185 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID vdd</lparam></gate>
<gate>
<ID>980</ID>
<type>DA_FROM</type>
<position>148.5,-164.5</position>
<input>
<ID>IN_0</ID>1186 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID gnd</lparam></gate>
<gate>
<ID>981</ID>
<type>DA_FROM</type>
<position>143.5,-168</position>
<input>
<ID>IN_0</ID>1187 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ldOut</lparam></gate>
<gate>
<ID>982</ID>
<type>DA_FROM</type>
<position>109,-9.5</position>
<input>
<ID>IN_0</ID>801 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID arBus</lparam></gate>
<gate>
<ID>983</ID>
<type>DA_FROM</type>
<position>109,-61.5</position>
<input>
<ID>IN_0</ID>1188 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID drBus</lparam></gate>
<gate>
<ID>984</ID>
<type>DA_FROM</type>
<position>109,-89.5</position>
<input>
<ID>IN_0</ID>755 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID acBus</lparam></gate>
<gate>
<ID>985</ID>
<type>DA_FROM</type>
<position>109.5,-121.5</position>
<input>
<ID>IN_0</ID>756 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID irBus</lparam></gate>
<gate>
<ID>986</ID>
<type>DA_FROM</type>
<position>153,-189.5</position>
<input>
<ID>IN_0</ID>754 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clrOut</lparam></gate>
<gate>
<ID>990</ID>
<type>AA_TOGGLE</type>
<position>40,0</position>
<output>
<ID>OUT_0</ID>1191 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>992</ID>
<type>BB_CLOCK</type>
<position>41,4.5</position>
<output>
<ID>CLK</ID>1192 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>994</ID>
<type>DE_TO</type>
<position>47,0</position>
<input>
<ID>IN_0</ID>1191 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID start</lparam></gate>
<gate>
<ID>995</ID>
<type>AA_LABEL</type>
<position>-34,11</position>
<gparam>LABEL_TEXT Datapath</gparam>
<gparam>TEXT_HEIGHT 10</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>758 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,6.5,108,6.5</points>
<connection>
<GID>819</GID>
<name>ADDRESS_2</name></connection>
<intersection>90 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>90,6.5,90,6.5</points>
<connection>
<GID>841</GID>
<name>IN_2</name></connection>
<intersection>6.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>837 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>107.5,-28.5,110.5,-28.5</points>
<connection>
<GID>855</GID>
<name>IN_2</name></connection>
<intersection>107.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>107.5,-29,107.5,-28.5</points>
<connection>
<GID>847</GID>
<name>OUT_2</name></connection>
<intersection>-28.5 0</intersection></vsegment></shape></wire>
<wire>
<ID>1144 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-108,63,-108</points>
<connection>
<GID>882</GID>
<name>IN_0</name></connection>
<connection>
<GID>857</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1165 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-173,69.5,-169.5</points>
<connection>
<GID>864</GID>
<name>clear</name></connection>
<intersection>-173 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-173,69.5,-173</points>
<connection>
<GID>898</GID>
<name>IN_0</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>832 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-51,104,-51</points>
<connection>
<GID>820</GID>
<name>OUT_3</name></connection>
<connection>
<GID>853</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1101 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-186,154,-186</points>
<connection>
<GID>836</GID>
<name>OUT_0</name></connection>
<connection>
<GID>875</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>768 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,9.5,108,9.5</points>
<connection>
<GID>819</GID>
<name>ADDRESS_5</name></connection>
<intersection>90 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>90,9.5,90,9.5</points>
<connection>
<GID>843</GID>
<name>IN_1</name></connection>
<intersection>9.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1117 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-176,164.5,-176</points>
<connection>
<GID>876</GID>
<name>IN_2</name></connection>
<connection>
<GID>878</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>767 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,15.5,108,15.5</points>
<connection>
<GID>819</GID>
<name>ADDRESS_11</name></connection>
<intersection>90 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>90,15.5,90,15.5</points>
<connection>
<GID>843</GID>
<name>IN_7</name></connection>
<intersection>15.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>840 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-25.5,108,-24.5</points>
<intersection>-25.5 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-25.5,110.5,-25.5</points>
<connection>
<GID>855</GID>
<name>IN_5</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-24.5,108,-24.5</points>
<connection>
<GID>845</GID>
<name>OUT_1</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>1173 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-41,69.5,-35.5</points>
<connection>
<GID>820</GID>
<name>count_up</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-35.5,69.5,-35.5</points>
<connection>
<GID>973</GID>
<name>IN_0</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1109 1110 1111 1112 1113 1114 1115 1116 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>158,-174.5,160.5,-174.5</points>
<connection>
<GID>874</GID>
<name>OUT</name></connection>
<connection>
<GID>878</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>776 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-23.5,73,-23.5</points>
<connection>
<GID>824</GID>
<name>OUT_6</name></connection>
<connection>
<GID>837</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>759 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,4.5,108,4.5</points>
<connection>
<GID>819</GID>
<name>ADDRESS_0</name></connection>
<intersection>90 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>90,4.5,90,4.5</points>
<connection>
<GID>841</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>757 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,5.5,108,5.5</points>
<connection>
<GID>819</GID>
<name>ADDRESS_1</name></connection>
<intersection>90 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>90,5.5,90,5.5</points>
<connection>
<GID>841</GID>
<name>IN_1</name></connection>
<intersection>5.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>761 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,14.5,108,14.5</points>
<connection>
<GID>819</GID>
<name>ADDRESS_10</name></connection>
<intersection>90 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>90,14.5,90,14.5</points>
<connection>
<GID>843</GID>
<name>IN_6</name></connection>
<intersection>14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>999 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-47,63.5,-47</points>
<connection>
<GID>848</GID>
<name>IN_7</name></connection>
<connection>
<GID>820</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>807 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-1,113.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_11</name></connection>
<intersection>-1 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-1,113.5,-1</points>
<intersection>113.5 0</intersection>
<intersection>113.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-1,113.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_11</name></connection>
<intersection>113.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>113.5,-1,113.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_11</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>1118 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-172,164.5,-172</points>
<connection>
<GID>876</GID>
<name>IN_6</name></connection>
<connection>
<GID>878</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>760 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,7.5,108,7.5</points>
<connection>
<GID>819</GID>
<name>ADDRESS_3</name></connection>
<intersection>90 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>90,7.5,90,7.5</points>
<connection>
<GID>841</GID>
<name>IN_3</name></connection>
<intersection>7.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>764 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,8.5,108,8.5</points>
<connection>
<GID>819</GID>
<name>ADDRESS_4</name></connection>
<intersection>90 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>90,8.5,90,8.5</points>
<connection>
<GID>843</GID>
<name>IN_0</name></connection>
<intersection>8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1176 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-62.5,67,-62</points>
<connection>
<GID>821</GID>
<name>load</name></connection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-62.5,67,-62.5</points>
<connection>
<GID>946</GID>
<name>IN_0</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>997 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-52,63.5,-52</points>
<connection>
<GID>848</GID>
<name>IN_2</name></connection>
<connection>
<GID>820</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>766 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,10.5,108,10.5</points>
<connection>
<GID>819</GID>
<name>ADDRESS_6</name></connection>
<intersection>90 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>90,10.5,90,10.5</points>
<connection>
<GID>843</GID>
<name>IN_2</name></connection>
<intersection>10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>993 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-50,63.5,-50</points>
<connection>
<GID>848</GID>
<name>IN_4</name></connection>
<connection>
<GID>820</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>762 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,11.5,108,11.5</points>
<connection>
<GID>819</GID>
<name>ADDRESS_7</name></connection>
<intersection>90 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>90,11.5,90,11.5</points>
<connection>
<GID>843</GID>
<name>IN_3</name></connection>
<intersection>11.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>765 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,12.5,108,12.5</points>
<connection>
<GID>819</GID>
<name>ADDRESS_8</name></connection>
<intersection>90 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>90,12.5,90,12.5</points>
<connection>
<GID>843</GID>
<name>IN_4</name></connection>
<intersection>12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>796 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-25.5,103.5,-25.5</points>
<connection>
<GID>849</GID>
<name>IN_0</name></connection>
<connection>
<GID>845</GID>
<name>IN_0</name></connection>
<intersection>98.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>98.5,-25.5,98.5,-15.5</points>
<connection>
<GID>905</GID>
<name>IN_0</name></connection>
<intersection>-25.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>763 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,13.5,108,13.5</points>
<connection>
<GID>819</GID>
<name>ADDRESS_9</name></connection>
<intersection>90 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>90,13.5,90,13.5</points>
<connection>
<GID>843</GID>
<name>IN_5</name></connection>
<intersection>13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>812 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-1,124.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_0</name></connection>
<intersection>-1 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,-1,124.5,-1</points>
<intersection>124.5 0</intersection>
<intersection>124.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,-1,124.5,-1</points>
<connection>
<GID>852</GID>
<name>Bus_in_0</name></connection>
<intersection>124.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>124.5,-1,124.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>1180 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-124,67.5,-122.5</points>
<connection>
<GID>861</GID>
<name>load</name></connection>
<intersection>-122.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-122.5,67.5,-122.5</points>
<connection>
<GID>966</GID>
<name>IN_0</name></connection>
<intersection>67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>817 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-1,123.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_1</name></connection>
<intersection>-1 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123.5,-1,123.5,-1</points>
<intersection>123.5 0</intersection>
<intersection>123.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-1,123.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_1</name></connection>
<intersection>123.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>123.5,-1,123.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>821 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-1,114.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_10</name></connection>
<intersection>-1 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-1,114.5,-1</points>
<intersection>114.5 0</intersection>
<intersection>114.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-1,114.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_10</name></connection>
<intersection>114.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114.5,-1,114.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_10</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>1000 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-45,63.5,-45</points>
<connection>
<GID>848</GID>
<name>IN_9</name></connection>
<connection>
<GID>820</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>808 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-1,112.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_12</name></connection>
<intersection>-1 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,-1,112.5,-1</points>
<intersection>112.5 0</intersection>
<intersection>112.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>112.5,-1,112.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_12</name></connection>
<intersection>112.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>112.5,-1,112.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_12</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>1146 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-106,63,-106</points>
<connection>
<GID>856</GID>
<name>IN_0</name></connection>
<connection>
<GID>857</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>811 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-1,111.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_13</name></connection>
<intersection>-1 2</intersection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,-1,111.5,-1</points>
<intersection>111.5 0</intersection>
<intersection>111.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-1,111.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_13</name></connection>
<intersection>111.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>111.5,-1,111.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_13</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>1149 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-100,63,-100</points>
<connection>
<GID>857</GID>
<name>IN_8</name></connection>
<connection>
<GID>885</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>816 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-1,110.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_14</name></connection>
<intersection>-1 2</intersection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110.5,-1,110.5,-1</points>
<intersection>110.5 0</intersection>
<intersection>110.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110.5,-1,110.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_14</name></connection>
<intersection>110.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110.5,-1,110.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_14</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>809 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-1,109.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_15</name></connection>
<intersection>-1 2</intersection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-1,109.5,-1</points>
<intersection>109.5 0</intersection>
<intersection>109.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,-1,109.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_15</name></connection>
<intersection>109.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>109.5,-1,109.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_15</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>1172 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-41,68.5,-38</points>
<connection>
<GID>820</GID>
<name>count_enable</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-38,68.5,-38</points>
<connection>
<GID>955</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1001 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-43,63.5,-43</points>
<connection>
<GID>848</GID>
<name>IN_11</name></connection>
<connection>
<GID>820</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>819 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-1,122.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_2</name></connection>
<intersection>-1 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-1,122.5,-1</points>
<intersection>122.5 0</intersection>
<intersection>122.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>122.5,-1,122.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_2</name></connection>
<intersection>122.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>122.5,-1,122.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>1026 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-69,63,-69</points>
<connection>
<GID>850</GID>
<name>IN_10</name></connection>
<connection>
<GID>821</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>813 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-1,121.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_3</name></connection>
<intersection>-1 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-1,121.5,-1</points>
<intersection>121.5 0</intersection>
<intersection>121.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121.5,-1,121.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_3</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>121.5,-1,121.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>1143 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,11.5,139.5,11.5</points>
<connection>
<GID>819</GID>
<name>write_clock</name></connection>
<intersection>135.5 3</intersection>
<intersection>139.5 36</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>135.5,-190.5,135.5,11.5</points>
<intersection>-190.5 31</intersection>
<intersection>-164 28</intersection>
<intersection>-144.5 27</intersection>
<intersection>-110.5 22</intersection>
<intersection>-80.5 17</intersection>
<intersection>-55.5 12</intersection>
<intersection>-32 8</intersection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>67,-32,135.5,-32</points>
<intersection>67 32</intersection>
<intersection>135.5 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>67.5,-55.5,135.5,-55.5</points>
<intersection>67.5 35</intersection>
<intersection>135.5 3</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>67,-80.5,135.5,-80.5</points>
<intersection>67 19</intersection>
<intersection>135.5 3</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>67,-81,67,-80.5</points>
<connection>
<GID>821</GID>
<name>clock</name></connection>
<intersection>-80.5 17</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>67,-110.5,135.5,-110.5</points>
<intersection>67 24</intersection>
<intersection>135.5 3</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>67,-110.5,67,-110</points>
<connection>
<GID>857</GID>
<name>clock</name></connection>
<intersection>-110.5 22</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>67.5,-144.5,135.5,-144.5</points>
<intersection>67.5 33</intersection>
<intersection>135.5 3</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>67.5,-164,135.5,-164</points>
<intersection>67.5 30</intersection>
<intersection>135.5 3</intersection></hsegment>
<vsegment>
<ID>30</ID>
<points>67.5,-169.5,67.5,-164</points>
<connection>
<GID>864</GID>
<name>clock</name></connection>
<intersection>-164 28</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>135.5,-190.5,147.5,-190.5</points>
<intersection>135.5 3</intersection>
<intersection>147.5 34</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>67,-32,67,-31.5</points>
<connection>
<GID>824</GID>
<name>clock</name></connection>
<intersection>-32 8</intersection></vsegment>
<vsegment>
<ID>33</ID>
<points>67.5,-144.5,67.5,-143</points>
<connection>
<GID>861</GID>
<name>clock</name></connection>
<intersection>-144.5 27</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>147.5,-190.5,147.5,-188</points>
<connection>
<GID>836</GID>
<name>clock</name></connection>
<intersection>-190.5 31</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>67.5,-56,67.5,-55.5</points>
<connection>
<GID>820</GID>
<name>clock</name></connection>
<intersection>-55.5 12</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>139.5,11.5,139.5,11.5</points>
<connection>
<GID>881</GID>
<name>IN_0</name></connection>
<intersection>11.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>814 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120.5,-1,120.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_4</name></connection>
<intersection>-1 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120.5,-1,120.5,-1</points>
<intersection>120.5 0</intersection>
<intersection>120.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120.5,-1,120.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_4</name></connection>
<intersection>120.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>120.5,-1,120.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_4</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>998 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-49,63.5,-49</points>
<connection>
<GID>848</GID>
<name>IN_5</name></connection>
<connection>
<GID>820</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>806 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-1,119.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_5</name></connection>
<intersection>-1 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,-1,119.5,-1</points>
<intersection>119.5 0</intersection>
<intersection>119.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119.5,-1,119.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_5</name></connection>
<intersection>119.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>119.5,-1,119.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_5</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>1161 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-57,69.5,-56</points>
<connection>
<GID>894</GID>
<name>IN_0</name></connection>
<connection>
<GID>820</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>820 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-1,118.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_6</name></connection>
<intersection>-1 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118.5,-1,118.5,-1</points>
<intersection>118.5 0</intersection>
<intersection>118.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>118.5,-1,118.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_6</name></connection>
<intersection>118.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>118.5,-1,118.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_6</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>810 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-1,117.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_7</name></connection>
<intersection>-1 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-1,117.5,-1</points>
<intersection>117.5 0</intersection>
<intersection>117.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>117.5,-1,117.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_7</name></connection>
<intersection>117.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>117.5,-1,117.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_7</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>815 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-1,116.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_8</name></connection>
<intersection>-1 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-1,116.5,-1</points>
<intersection>116.5 0</intersection>
<intersection>116.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116.5,-1,116.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_8</name></connection>
<intersection>116.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116.5,-1,116.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_8</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>818 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-1,115.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_IN_9</name></connection>
<intersection>-1 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-1,115.5,-1</points>
<intersection>115.5 0</intersection>
<intersection>115.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115.5,-1,115.5,-1</points>
<connection>
<GID>852</GID>
<name>IN_9</name></connection>
<intersection>115.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>115.5,-1,115.5,-1</points>
<connection>
<GID>819</GID>
<name>DATA_OUT_9</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>1167 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,7.5,138.5,9.5</points>
<intersection>7.5 2</intersection>
<intersection>9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,9.5,138.5,9.5</points>
<connection>
<GID>819</GID>
<name>ENABLE_0</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138.5,7.5,139.5,7.5</points>
<connection>
<GID>900</GID>
<name>IN_0</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1166 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,10.5,139.5,10.5</points>
<connection>
<GID>819</GID>
<name>write_enable</name></connection>
<intersection>139.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>139.5,9.5,139.5,10.5</points>
<connection>
<GID>899</GID>
<name>IN_0</name></connection>
<intersection>10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1145 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-107,63,-107</points>
<connection>
<GID>857</GID>
<name>IN_1</name></connection>
<connection>
<GID>830</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>996 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-54,63.5,-54</points>
<connection>
<GID>848</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>820</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>992 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-53,63.5,-53</points>
<connection>
<GID>848</GID>
<name>IN_1</name></connection>
<connection>
<GID>820</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>991 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-44,63.5,-44</points>
<connection>
<GID>848</GID>
<name>IN_10</name></connection>
<connection>
<GID>820</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>995 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-51,63.5,-51</points>
<connection>
<GID>848</GID>
<name>IN_3</name></connection>
<connection>
<GID>820</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>990 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-48,63.5,-48</points>
<connection>
<GID>848</GID>
<name>IN_6</name></connection>
<connection>
<GID>820</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>994 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-46,63.5,-46</points>
<connection>
<GID>848</GID>
<name>IN_8</name></connection>
<connection>
<GID>820</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1171 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-41,67.5,-40</points>
<connection>
<GID>820</GID>
<name>load</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-40,67.5,-40</points>
<connection>
<GID>972</GID>
<name>IN_0</name></connection>
<intersection>67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>833 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-54,104,-54</points>
<connection>
<GID>820</GID>
<name>OUT_0</name></connection>
<connection>
<GID>853</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1139 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-173,179,-173</points>
<connection>
<GID>877</GID>
<name>IN_5</name></connection>
<connection>
<GID>879</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>834 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-53,104,-53</points>
<connection>
<GID>820</GID>
<name>OUT_1</name></connection>
<connection>
<GID>853</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1034 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-132,63.5,-132</points>
<connection>
<GID>870</GID>
<name>IN_9</name></connection>
<connection>
<GID>861</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>827 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-44,104,-44</points>
<connection>
<GID>820</GID>
<name>OUT_10</name></connection>
<connection>
<GID>854</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>830 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-43,104,-43</points>
<connection>
<GID>820</GID>
<name>OUT_11</name></connection>
<connection>
<GID>854</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>831 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-52,104,-52</points>
<connection>
<GID>820</GID>
<name>OUT_2</name></connection>
<connection>
<GID>853</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1029 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-140,63.5,-140</points>
<connection>
<GID>870</GID>
<name>IN_1</name></connection>
<connection>
<GID>861</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>824 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-50,104,-50</points>
<connection>
<GID>820</GID>
<name>OUT_4</name></connection>
<connection>
<GID>854</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1015 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-79,63,-79</points>
<connection>
<GID>850</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>821</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>823 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-49,104,-49</points>
<connection>
<GID>820</GID>
<name>OUT_5</name></connection>
<connection>
<GID>854</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1017 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-67,63,-67</points>
<connection>
<GID>850</GID>
<name>IN_12</name></connection>
<connection>
<GID>821</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1188 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-62.5,106,-61.5</points>
<connection>
<GID>831</GID>
<name>ENABLE_0</name></connection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-61.5,107,-61.5</points>
<connection>
<GID>983</GID>
<name>IN_0</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>825 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-48,104,-48</points>
<connection>
<GID>820</GID>
<name>OUT_6</name></connection>
<connection>
<GID>854</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>826 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-47,104,-47</points>
<connection>
<GID>820</GID>
<name>OUT_7</name></connection>
<connection>
<GID>854</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>829 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-46,104,-46</points>
<connection>
<GID>820</GID>
<name>OUT_8</name></connection>
<connection>
<GID>854</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1041 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-128,63.5,-128</points>
<connection>
<GID>870</GID>
<name>IN_13</name></connection>
<connection>
<GID>861</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1020 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-68,63,-68</points>
<connection>
<GID>850</GID>
<name>IN_11</name></connection>
<connection>
<GID>821</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>828 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-45,104,-45</points>
<connection>
<GID>820</GID>
<name>OUT_9</name></connection>
<connection>
<GID>854</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>845 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-20.5,109.5,-19.5</points>
<intersection>-20.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-19.5,109.5,-19.5</points>
<connection>
<GID>845</GID>
<name>OUT_6</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,-20.5,110.5,-20.5</points>
<connection>
<GID>855</GID>
<name>IN_10</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1024 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-78,63,-78</points>
<connection>
<GID>850</GID>
<name>IN_1</name></connection>
<connection>
<GID>821</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1018 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-66,63,-66</points>
<connection>
<GID>850</GID>
<name>IN_13</name></connection>
<connection>
<GID>821</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1019 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-65,63,-65</points>
<connection>
<GID>850</GID>
<name>IN_14</name></connection>
<connection>
<GID>821</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1028 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-64,63,-64</points>
<connection>
<GID>850</GID>
<name>IN_15</name></connection>
<connection>
<GID>821</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1023 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-77,63,-77</points>
<connection>
<GID>850</GID>
<name>IN_2</name></connection>
<connection>
<GID>821</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1022 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-76,63,-76</points>
<connection>
<GID>850</GID>
<name>IN_3</name></connection>
<connection>
<GID>821</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>850 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-50,111,-50</points>
<connection>
<GID>854</GID>
<name>OUT_0</name></connection>
<connection>
<GID>827</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1027 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-75,63,-75</points>
<connection>
<GID>850</GID>
<name>IN_4</name></connection>
<connection>
<GID>821</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1014 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-74,63,-74</points>
<connection>
<GID>850</GID>
<name>IN_5</name></connection>
<connection>
<GID>821</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1021 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-73,63,-73</points>
<connection>
<GID>850</GID>
<name>IN_6</name></connection>
<connection>
<GID>821</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1192 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,4.5,45,4.5</points>
<connection>
<GID>868</GID>
<name>IN_0</name></connection>
<connection>
<GID>992</GID>
<name>CLK</name></connection></vsegment></shape></wire>
<wire>
<ID>1013 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-72,63,-72</points>
<connection>
<GID>850</GID>
<name>IN_7</name></connection>
<connection>
<GID>821</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1016 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-71,63,-71</points>
<connection>
<GID>850</GID>
<name>IN_8</name></connection>
<connection>
<GID>821</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1004 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-21.5,63,-21.5</points>
<connection>
<GID>846</GID>
<name>IN_8</name></connection>
<connection>
<GID>824</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1025 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-70,63,-70</points>
<connection>
<GID>850</GID>
<name>IN_9</name></connection>
<connection>
<GID>821</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>955 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-155.5,104,-155.5</points>
<connection>
<GID>864</GID>
<name>OUT_12</name></connection>
<connection>
<GID>866</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1162 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-82.5,69,-81</points>
<connection>
<GID>821</GID>
<name>clear</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-82.5,69,-82.5</points>
<connection>
<GID>895</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>1175 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-62,68,-60.5</points>
<connection>
<GID>821</GID>
<name>count_enable</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-60.5,68,-60.5</points>
<connection>
<GID>974</GID>
<name>IN_0</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>1174 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-62,69,-58.5</points>
<connection>
<GID>821</GID>
<name>count_up</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-58.5,69,-58.5</points>
<connection>
<GID>940</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>867 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-79,104,-79</points>
<connection>
<GID>821</GID>
<name>OUT_0</name></connection>
<connection>
<GID>831</GID>
<name>IN_0</name></connection>
<intersection>103.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>103.5,-79,103.5,-63.5</points>
<connection>
<GID>913</GID>
<name>IN_0</name></connection>
<intersection>-79 1</intersection></vsegment></shape></wire>
<wire>
<ID>871 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-78,104,-78</points>
<connection>
<GID>821</GID>
<name>OUT_1</name></connection>
<connection>
<GID>831</GID>
<name>IN_1</name></connection>
<intersection>101.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>101.5,-78,101.5,-63.5</points>
<connection>
<GID>914</GID>
<name>IN_0</name></connection>
<intersection>-78 1</intersection></vsegment></shape></wire>
<wire>
<ID>864 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-69,104,-69</points>
<connection>
<GID>821</GID>
<name>OUT_10</name></connection>
<connection>
<GID>831</GID>
<name>IN_10</name></connection>
<intersection>83.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>83.5,-69,83.5,-63.5</points>
<connection>
<GID>923</GID>
<name>IN_0</name></connection>
<intersection>-69 1</intersection></vsegment></shape></wire>
<wire>
<ID>870 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-68,104,-68</points>
<connection>
<GID>821</GID>
<name>OUT_11</name></connection>
<connection>
<GID>831</GID>
<name>IN_11</name></connection>
<intersection>81.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>81.5,-68,81.5,-63.5</points>
<connection>
<GID>924</GID>
<name>IN_0</name></connection>
<intersection>-68 1</intersection></vsegment></shape></wire>
<wire>
<ID>859 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-67,104,-67</points>
<connection>
<GID>821</GID>
<name>OUT_12</name></connection>
<connection>
<GID>831</GID>
<name>IN_12</name></connection>
<intersection>79.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>79.5,-67,79.5,-63.5</points>
<connection>
<GID>925</GID>
<name>IN_0</name></connection>
<intersection>-67 1</intersection></vsegment></shape></wire>
<wire>
<ID>860 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-66,104,-66</points>
<connection>
<GID>821</GID>
<name>OUT_13</name></connection>
<connection>
<GID>831</GID>
<name>IN_13</name></connection>
<intersection>77.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>77.5,-66,77.5,-63.5</points>
<connection>
<GID>926</GID>
<name>IN_0</name></connection>
<intersection>-66 1</intersection></vsegment></shape></wire>
<wire>
<ID>873 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-65,104,-65</points>
<connection>
<GID>821</GID>
<name>OUT_14</name></connection>
<connection>
<GID>831</GID>
<name>IN_14</name></connection>
<intersection>75.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>75.5,-65,75.5,-63.5</points>
<connection>
<GID>927</GID>
<name>IN_0</name></connection>
<intersection>-65 1</intersection></vsegment></shape></wire>
<wire>
<ID>1051 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-164.5,63.5,-164.5</points>
<connection>
<GID>871</GID>
<name>IN_3</name></connection>
<connection>
<GID>864</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>874 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-64,104,-64</points>
<connection>
<GID>821</GID>
<name>OUT_15</name></connection>
<connection>
<GID>831</GID>
<name>IN_15</name></connection>
<intersection>73.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>73.5,-64,73.5,-63.5</points>
<connection>
<GID>928</GID>
<name>IN_0</name></connection>
<intersection>-64 1</intersection></vsegment></shape></wire>
<wire>
<ID>865 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-77,104,-77</points>
<connection>
<GID>821</GID>
<name>OUT_2</name></connection>
<connection>
<GID>831</GID>
<name>IN_2</name></connection>
<intersection>99.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>99.5,-77,99.5,-63.5</points>
<connection>
<GID>915</GID>
<name>IN_0</name></connection>
<intersection>-77 1</intersection></vsegment></shape></wire>
<wire>
<ID>1043 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-130,63.5,-130</points>
<connection>
<GID>870</GID>
<name>IN_11</name></connection>
<connection>
<GID>861</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>866 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-76,104,-76</points>
<connection>
<GID>821</GID>
<name>OUT_3</name></connection>
<connection>
<GID>831</GID>
<name>IN_3</name></connection>
<intersection>97.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>97.5,-76,97.5,-63.5</points>
<connection>
<GID>916</GID>
<name>IN_0</name></connection>
<intersection>-76 1</intersection></vsegment></shape></wire>
<wire>
<ID>868 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-75,104,-75</points>
<connection>
<GID>821</GID>
<name>OUT_4</name></connection>
<connection>
<GID>831</GID>
<name>IN_4</name></connection>
<intersection>95.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>95.5,-75,95.5,-63.5</points>
<connection>
<GID>917</GID>
<name>IN_0</name></connection>
<intersection>-75 1</intersection></vsegment></shape></wire>
<wire>
<ID>862 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-74,104,-74</points>
<connection>
<GID>821</GID>
<name>OUT_5</name></connection>
<connection>
<GID>831</GID>
<name>IN_5</name></connection>
<intersection>93.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>93.5,-74,93.5,-63.5</points>
<connection>
<GID>918</GID>
<name>IN_0</name></connection>
<intersection>-74 1</intersection></vsegment></shape></wire>
<wire>
<ID>1048 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-157.5,63.5,-157.5</points>
<connection>
<GID>871</GID>
<name>IN_10</name></connection>
<connection>
<GID>864</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>869 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-73,104,-73</points>
<connection>
<GID>821</GID>
<name>OUT_6</name></connection>
<connection>
<GID>831</GID>
<name>IN_6</name></connection>
<intersection>91.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>91.5,-73,91.5,-63.5</points>
<connection>
<GID>919</GID>
<name>IN_0</name></connection>
<intersection>-73 1</intersection></vsegment></shape></wire>
<wire>
<ID>872 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-72,104,-72</points>
<connection>
<GID>821</GID>
<name>OUT_7</name></connection>
<connection>
<GID>831</GID>
<name>IN_7</name></connection>
<intersection>89.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>89.5,-72,89.5,-63.5</points>
<connection>
<GID>920</GID>
<name>IN_0</name></connection>
<intersection>-72 1</intersection></vsegment></shape></wire>
<wire>
<ID>863 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-71,104,-71</points>
<connection>
<GID>821</GID>
<name>OUT_8</name></connection>
<connection>
<GID>831</GID>
<name>IN_8</name></connection>
<intersection>87.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>87.5,-71,87.5,-63.5</points>
<connection>
<GID>921</GID>
<name>IN_0</name></connection>
<intersection>-71 1</intersection></vsegment></shape></wire>
<wire>
<ID>1040 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-126,63.5,-126</points>
<connection>
<GID>870</GID>
<name>IN_15</name></connection>
<connection>
<GID>861</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>861 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-70,104,-70</points>
<connection>
<GID>821</GID>
<name>OUT_9</name></connection>
<connection>
<GID>831</GID>
<name>IN_9</name></connection>
<intersection>85.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>85.5,-70,85.5,-63.5</points>
<connection>
<GID>922</GID>
<name>IN_0</name></connection>
<intersection>-70 1</intersection></vsegment></shape></wire>
<wire>
<ID>1179 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-91,69,-86.5</points>
<connection>
<GID>857</GID>
<name>count_up</name></connection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-86.5,69,-86.5</points>
<connection>
<GID>976</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>1002 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-29.5,63,-29.5</points>
<connection>
<GID>846</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>824</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1184 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-150.5,68.5,-148</points>
<connection>
<GID>864</GID>
<name>count_enable</name></connection>
<intersection>-148 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-148,68.5,-148</points>
<connection>
<GID>949</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1005 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-28.5,63,-28.5</points>
<connection>
<GID>846</GID>
<name>IN_1</name></connection>
<connection>
<GID>824</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1033 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-139,63.5,-139</points>
<connection>
<GID>870</GID>
<name>IN_2</name></connection>
<connection>
<GID>861</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1012 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-19.5,63,-19.5</points>
<connection>
<GID>846</GID>
<name>IN_10</name></connection>
<connection>
<GID>824</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1011 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-18.5,63,-18.5</points>
<connection>
<GID>846</GID>
<name>IN_11</name></connection>
<connection>
<GID>824</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1008 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-27.5,63,-27.5</points>
<connection>
<GID>846</GID>
<name>IN_2</name></connection>
<connection>
<GID>824</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1006 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-26.5,63,-26.5</points>
<connection>
<GID>846</GID>
<name>IN_3</name></connection>
<connection>
<GID>824</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1009 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-25.5,63,-25.5</points>
<connection>
<GID>846</GID>
<name>IN_4</name></connection>
<connection>
<GID>824</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1187 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,-169,147.5,-168</points>
<connection>
<GID>836</GID>
<name>load</name></connection>
<intersection>-168 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,-168,147.5,-168</points>
<connection>
<GID>981</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1010 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-24.5,63,-24.5</points>
<connection>
<GID>846</GID>
<name>IN_5</name></connection>
<connection>
<GID>824</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1007 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-23.5,63,-23.5</points>
<connection>
<GID>846</GID>
<name>IN_6</name></connection>
<connection>
<GID>824</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1003 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-22.5,63,-22.5</points>
<connection>
<GID>846</GID>
<name>IN_7</name></connection>
<connection>
<GID>824</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1190 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-20.5,63,-20.5</points>
<connection>
<GID>846</GID>
<name>IN_9</name></connection>
<connection>
<GID>824</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>981 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-158.5,111,-158.5</points>
<connection>
<GID>866</GID>
<name>OUT_9</name></connection>
<connection>
<GID>865</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1160 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>66.5,-32.5,69,-32.5</points>
<connection>
<GID>893</GID>
<name>IN_0</name></connection>
<intersection>69 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>69,-32.5,69,-31.5</points>
<connection>
<GID>824</GID>
<name>clear</name></connection>
<intersection>-32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1169 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-16.5,68,-13.5</points>
<connection>
<GID>824</GID>
<name>count_enable</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-13.5,68,-13.5</points>
<connection>
<GID>970</GID>
<name>IN_0</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>835 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>107.5,-30.5,110.5,-30.5</points>
<connection>
<GID>855</GID>
<name>Bus_in_0</name></connection>
<intersection>107.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>107.5,-31,107.5,-30.5</points>
<connection>
<GID>847</GID>
<name>OUT_0</name></connection>
<intersection>-30.5 0</intersection></vsegment></shape></wire>
<wire>
<ID>1170 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-16.5,69,-11.5</points>
<connection>
<GID>824</GID>
<name>count_up</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-11.5,69,-11.5</points>
<connection>
<GID>971</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>989 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,10.5,44,10.5</points>
<connection>
<GID>844</GID>
<name>IN_0</name></connection>
<intersection>40 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>40,10,40,10.5</points>
<connection>
<GID>842</GID>
<name>OUT_0</name></connection>
<intersection>10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1168 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>66.5,-15.5,67,-15.5</points>
<connection>
<GID>969</GID>
<name>IN_0</name></connection>
<intersection>67 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>67,-16.5,67,-15.5</points>
<connection>
<GID>824</GID>
<name>load</name></connection>
<intersection>-15.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>777 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-29.5,73,-29.5</points>
<connection>
<GID>824</GID>
<name>OUT_0</name></connection>
<connection>
<GID>839</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>779 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-28.5,73,-28.5</points>
<connection>
<GID>824</GID>
<name>OUT_1</name></connection>
<connection>
<GID>839</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>775 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-19.5,73,-19.5</points>
<connection>
<GID>824</GID>
<name>OUT_10</name></connection>
<connection>
<GID>837</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>1106 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-181,154,-181</points>
<connection>
<GID>836</GID>
<name>OUT_5</name></connection>
<connection>
<GID>875</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>771 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-18.5,73,-18.5</points>
<connection>
<GID>824</GID>
<name>OUT_11</name></connection>
<connection>
<GID>837</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>778 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-27.5,73,-27.5</points>
<connection>
<GID>824</GID>
<name>OUT_2</name></connection>
<connection>
<GID>839</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>780 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-26.5,73,-26.5</points>
<connection>
<GID>824</GID>
<name>OUT_3</name></connection>
<connection>
<GID>839</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>773 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-25.5,73,-25.5</points>
<connection>
<GID>824</GID>
<name>OUT_4</name></connection>
<connection>
<GID>837</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>772 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-24.5,73,-24.5</points>
<connection>
<GID>824</GID>
<name>OUT_5</name></connection>
<connection>
<GID>837</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1075 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-174,143.5,-174</points>
<connection>
<GID>836</GID>
<name>IN_12</name></connection>
<connection>
<GID>872</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>770 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-22.5,73,-22.5</points>
<connection>
<GID>824</GID>
<name>OUT_7</name></connection>
<connection>
<GID>837</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>769 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-21.5,73,-21.5</points>
<connection>
<GID>824</GID>
<name>OUT_8</name></connection>
<connection>
<GID>837</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>774 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-20.5,73,-20.5</points>
<connection>
<GID>824</GID>
<name>OUT_9</name></connection>
<connection>
<GID>837</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>1035 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-141,63.5,-141</points>
<connection>
<GID>870</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>861</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>858 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-54,111,-54</points>
<connection>
<GID>853</GID>
<name>OUT_0</name></connection>
<connection>
<GID>827</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1189 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-151,106,-150</points>
<connection>
<GID>866</GID>
<name>ENABLE_0</name></connection>
<intersection>-150 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-150,106,-150</points>
<connection>
<GID>873</GID>
<name>IN_0</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>856 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-53,111,-53</points>
<connection>
<GID>853</GID>
<name>OUT_1</name></connection>
<connection>
<GID>827</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>849 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-44,111,-44</points>
<connection>
<GID>854</GID>
<name>OUT_6</name></connection>
<connection>
<GID>827</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>847 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-43,111,-43</points>
<connection>
<GID>854</GID>
<name>OUT_7</name></connection>
<connection>
<GID>827</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>857 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-52,111,-52</points>
<connection>
<GID>853</GID>
<name>OUT_2</name></connection>
<connection>
<GID>827</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>855 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-51,111,-51</points>
<connection>
<GID>853</GID>
<name>OUT_3</name></connection>
<connection>
<GID>827</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1032 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-133,63.5,-133</points>
<connection>
<GID>870</GID>
<name>IN_8</name></connection>
<connection>
<GID>861</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>853 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-49,111,-49</points>
<connection>
<GID>854</GID>
<name>OUT_1</name></connection>
<connection>
<GID>827</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1186 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-169,148.5,-166.5</points>
<connection>
<GID>836</GID>
<name>count_enable</name></connection>
<connection>
<GID>980</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>851 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-48,111,-48</points>
<connection>
<GID>854</GID>
<name>OUT_2</name></connection>
<connection>
<GID>827</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>854 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-47,111,-47</points>
<connection>
<GID>854</GID>
<name>OUT_3</name></connection>
<connection>
<GID>827</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>852 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-46,111,-46</points>
<connection>
<GID>854</GID>
<name>OUT_4</name></connection>
<connection>
<GID>827</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1181 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-124,68.5,-120.5</points>
<connection>
<GID>861</GID>
<name>count_enable</name></connection>
<intersection>-120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-120.5,68.5,-120.5</points>
<connection>
<GID>977</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>848 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-45,111,-45</points>
<connection>
<GID>854</GID>
<name>OUT_5</name></connection>
<connection>
<GID>827</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117,-178.5,117,-5</points>
<connection>
<GID>852</GID>
<name>OUT</name></connection>
<intersection>-178.5 11</intersection>
<intersection>-160 16</intersection>
<intersection>-133.5 9</intersection>
<intersection>-100.5 7</intersection>
<intersection>-71.5 5</intersection>
<intersection>-46.5 3</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-23,117,-23</points>
<connection>
<GID>855</GID>
<name>OUT</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>115,-46.5,117,-46.5</points>
<connection>
<GID>827</GID>
<name>OUT</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>114.5,-71.5,117,-71.5</points>
<connection>
<GID>829</GID>
<name>OUT</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>114.5,-100.5,117,-100.5</points>
<connection>
<GID>834</GID>
<name>OUT</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>115,-133.5,117,-133.5</points>
<connection>
<GID>862</GID>
<name>OUT</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>41,-178.5,137.5,-178.5</points>
<connection>
<GID>872</GID>
<name>OUT</name></connection>
<intersection>41 14</intersection>
<intersection>117 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>41,-178.5,41,-22</points>
<intersection>-178.5 11</intersection>
<intersection>-160 17</intersection>
<intersection>-133.5 19</intersection>
<intersection>-71.5 23</intersection>
<intersection>-46.5 25</intersection>
<intersection>-22 27</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>115,-160,117,-160</points>
<connection>
<GID>865</GID>
<name>OUT</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>41,-160,55.5,-160</points>
<connection>
<GID>871</GID>
<name>OUT</name></connection>
<intersection>41 14</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>41,-133.5,55.5,-133.5</points>
<connection>
<GID>870</GID>
<name>OUT</name></connection>
<intersection>41 14</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>41,-71.5,54.5,-71.5</points>
<connection>
<GID>850</GID>
<name>OUT</name></connection>
<intersection>41 14</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>41,-46.5,54.5,-46.5</points>
<connection>
<GID>848</GID>
<name>OUT</name></connection>
<intersection>41 14</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>41,-22,54,-22</points>
<connection>
<GID>846</GID>
<name>OUT</name></connection>
<intersection>41 14</intersection></hsegment></shape></wire>
<wire>
<ID>932 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-137,105.5,-137</points>
<connection>
<GID>861</GID>
<name>OUT_4</name></connection>
<connection>
<GID>863</GID>
<name>IN_4</name></connection>
<intersection>96.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>96.5,-137,96.5,-124.5</points>
<connection>
<GID>953</GID>
<name>IN_0</name></connection>
<intersection>-137 1</intersection></vsegment></shape></wire>
<wire>
<ID>967 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-166.5,104,-166.5</points>
<connection>
<GID>864</GID>
<name>OUT_1</name></connection>
<connection>
<GID>866</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>909 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-101,110.5,-101</points>
<connection>
<GID>859</GID>
<name>OUT_7</name></connection>
<connection>
<GID>834</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>883 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-68,110.5,-68</points>
<connection>
<GID>831</GID>
<name>OUT_11</name></connection>
<connection>
<GID>829</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>914 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-107,110.5,-107</points>
<connection>
<GID>859</GID>
<name>OUT_1</name></connection>
<connection>
<GID>834</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1067 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-186,143.5,-186</points>
<connection>
<GID>836</GID>
<name>IN_0</name></connection>
<connection>
<GID>872</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>890 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-79,110.5,-79</points>
<connection>
<GID>831</GID>
<name>OUT_0</name></connection>
<connection>
<GID>829</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1059 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-153.5,63.5,-153.5</points>
<connection>
<GID>871</GID>
<name>IN_14</name></connection>
<connection>
<GID>864</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>882 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-78,110.5,-78</points>
<connection>
<GID>831</GID>
<name>OUT_1</name></connection>
<connection>
<GID>829</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>881 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-69,110.5,-69</points>
<connection>
<GID>831</GID>
<name>OUT_10</name></connection>
<connection>
<GID>829</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>884 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-67,110.5,-67</points>
<connection>
<GID>831</GID>
<name>OUT_12</name></connection>
<connection>
<GID>829</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>879 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-66,110.5,-66</points>
<connection>
<GID>831</GID>
<name>OUT_13</name></connection>
<connection>
<GID>829</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>887 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-65,110.5,-65</points>
<connection>
<GID>831</GID>
<name>OUT_14</name></connection>
<connection>
<GID>829</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>886 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-64,110.5,-64</points>
<connection>
<GID>831</GID>
<name>OUT_15</name></connection>
<connection>
<GID>829</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1093 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-172,154,-172</points>
<connection>
<GID>836</GID>
<name>OUT_14</name></connection>
<connection>
<GID>874</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>888 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-77,110.5,-77</points>
<connection>
<GID>831</GID>
<name>OUT_2</name></connection>
<connection>
<GID>829</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>880 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-76,110.5,-76</points>
<connection>
<GID>831</GID>
<name>OUT_3</name></connection>
<connection>
<GID>829</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>876 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-75,110.5,-75</points>
<connection>
<GID>831</GID>
<name>OUT_4</name></connection>
<connection>
<GID>829</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>875 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-74,110.5,-74</points>
<connection>
<GID>831</GID>
<name>OUT_5</name></connection>
<connection>
<GID>829</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>878 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-73,110.5,-73</points>
<connection>
<GID>831</GID>
<name>OUT_6</name></connection>
<connection>
<GID>829</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1056 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-166.5,63.5,-166.5</points>
<connection>
<GID>871</GID>
<name>IN_1</name></connection>
<connection>
<GID>864</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>877 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-72,110.5,-72</points>
<connection>
<GID>831</GID>
<name>OUT_7</name></connection>
<connection>
<GID>829</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>889 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-71,110.5,-71</points>
<connection>
<GID>831</GID>
<name>OUT_8</name></connection>
<connection>
<GID>829</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1064 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-171,143.5,-171</points>
<connection>
<GID>836</GID>
<name>IN_15</name></connection>
<connection>
<GID>872</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>885 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-70,110.5,-70</points>
<connection>
<GID>831</GID>
<name>OUT_9</name></connection>
<connection>
<GID>829</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1159 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-105,63,-105</points>
<connection>
<GID>857</GID>
<name>IN_3</name></connection>
<connection>
<GID>833</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1099 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-176,154,-176</points>
<connection>
<GID>836</GID>
<name>OUT_10</name></connection>
<connection>
<GID>874</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>922 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-108,110.5,-108</points>
<connection>
<GID>859</GID>
<name>OUT_0</name></connection>
<connection>
<GID>834</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>913 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-98,110.5,-98</points>
<connection>
<GID>859</GID>
<name>OUT_10</name></connection>
<connection>
<GID>834</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>915 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-97,110.5,-97</points>
<connection>
<GID>859</GID>
<name>OUT_11</name></connection>
<connection>
<GID>834</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1065 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-177,143.5,-177</points>
<connection>
<GID>836</GID>
<name>IN_9</name></connection>
<connection>
<GID>872</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>916 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-96,110.5,-96</points>
<connection>
<GID>859</GID>
<name>OUT_12</name></connection>
<connection>
<GID>834</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>911 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-95,110.5,-95</points>
<connection>
<GID>859</GID>
<name>OUT_13</name></connection>
<connection>
<GID>834</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>919 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-94,110.5,-94</points>
<connection>
<GID>859</GID>
<name>OUT_14</name></connection>
<connection>
<GID>834</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>918 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-93,110.5,-93</points>
<connection>
<GID>859</GID>
<name>OUT_15</name></connection>
<connection>
<GID>834</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>920 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-106,110.5,-106</points>
<connection>
<GID>859</GID>
<name>OUT_2</name></connection>
<connection>
<GID>834</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>912 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-105,110.5,-105</points>
<connection>
<GID>859</GID>
<name>OUT_3</name></connection>
<connection>
<GID>834</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1057 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-162.5,63.5,-162.5</points>
<connection>
<GID>871</GID>
<name>IN_5</name></connection>
<connection>
<GID>864</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>908 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-104,110.5,-104</points>
<connection>
<GID>859</GID>
<name>OUT_4</name></connection>
<connection>
<GID>834</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>907 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-103,110.5,-103</points>
<connection>
<GID>859</GID>
<name>OUT_5</name></connection>
<connection>
<GID>834</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>910 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-102,110.5,-102</points>
<connection>
<GID>859</GID>
<name>OUT_6</name></connection>
<connection>
<GID>834</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>921 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-100,110.5,-100</points>
<connection>
<GID>859</GID>
<name>OUT_8</name></connection>
<connection>
<GID>834</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1096 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-174,154,-174</points>
<connection>
<GID>836</GID>
<name>OUT_12</name></connection>
<connection>
<GID>874</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>917 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-99,110.5,-99</points>
<connection>
<GID>859</GID>
<name>OUT_9</name></connection>
<connection>
<GID>834</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1066 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-185,143.5,-185</points>
<connection>
<GID>836</GID>
<name>IN_1</name></connection>
<connection>
<GID>872</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1063 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-176,143.5,-176</points>
<connection>
<GID>836</GID>
<name>IN_10</name></connection>
<connection>
<GID>872</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>924 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-128,105.5,-128</points>
<connection>
<GID>861</GID>
<name>OUT_13</name></connection>
<connection>
<GID>863</GID>
<name>IN_13</name></connection>
<intersection>78.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>78.5,-128,78.5,-124.5</points>
<connection>
<GID>965</GID>
<name>IN_0</name></connection>
<intersection>-128 1</intersection></vsegment></shape></wire>
<wire>
<ID>1073 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-175,143.5,-175</points>
<connection>
<GID>836</GID>
<name>IN_11</name></connection>
<connection>
<GID>872</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>893 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-99,105,-99</points>
<connection>
<GID>857</GID>
<name>OUT_9</name></connection>
<connection>
<GID>859</GID>
<name>IN_9</name></connection>
<intersection>86 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>86,-99,86,-91</points>
<connection>
<GID>938</GID>
<name>IN_0</name></connection>
<intersection>-99 1</intersection></vsegment></shape></wire>
<wire>
<ID>1072 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-173,143.5,-173</points>
<connection>
<GID>836</GID>
<name>IN_13</name></connection>
<connection>
<GID>872</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1076 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-172,143.5,-172</points>
<connection>
<GID>836</GID>
<name>IN_14</name></connection>
<connection>
<GID>872</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1074 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-184,143.5,-184</points>
<connection>
<GID>836</GID>
<name>IN_2</name></connection>
<connection>
<GID>872</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1068 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-183,143.5,-183</points>
<connection>
<GID>836</GID>
<name>IN_3</name></connection>
<connection>
<GID>872</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1061 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-182,143.5,-182</points>
<connection>
<GID>836</GID>
<name>IN_4</name></connection>
<connection>
<GID>872</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1062 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-181,143.5,-181</points>
<connection>
<GID>836</GID>
<name>IN_5</name></connection>
<connection>
<GID>872</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1069 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-180,143.5,-180</points>
<connection>
<GID>836</GID>
<name>IN_6</name></connection>
<connection>
<GID>872</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1070 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-179,143.5,-179</points>
<connection>
<GID>836</GID>
<name>IN_7</name></connection>
<connection>
<GID>872</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1071 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-178,143.5,-178</points>
<connection>
<GID>836</GID>
<name>IN_8</name></connection>
<connection>
<GID>872</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>754 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,-189.5,149.5,-188</points>
<connection>
<GID>836</GID>
<name>clear</name></connection>
<intersection>-189.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149.5,-189.5,151,-189.5</points>
<connection>
<GID>986</GID>
<name>IN_0</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1102 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-185,154,-185</points>
<connection>
<GID>836</GID>
<name>OUT_1</name></connection>
<connection>
<GID>875</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1100 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-175,154,-175</points>
<connection>
<GID>836</GID>
<name>OUT_11</name></connection>
<connection>
<GID>874</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1094 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-173,154,-173</points>
<connection>
<GID>836</GID>
<name>OUT_13</name></connection>
<connection>
<GID>874</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1097 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-171,154,-171</points>
<connection>
<GID>836</GID>
<name>OUT_15</name></connection>
<connection>
<GID>874</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1103 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-184,154,-184</points>
<connection>
<GID>836</GID>
<name>OUT_2</name></connection>
<connection>
<GID>875</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1105 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-183,154,-183</points>
<connection>
<GID>836</GID>
<name>OUT_3</name></connection>
<connection>
<GID>875</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>925 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-132,105.5,-132</points>
<connection>
<GID>861</GID>
<name>OUT_9</name></connection>
<connection>
<GID>863</GID>
<name>IN_9</name></connection>
<intersection>86.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>86.5,-132,86.5,-124.5</points>
<connection>
<GID>960</GID>
<name>IN_0</name></connection>
<intersection>-132 1</intersection></vsegment></shape></wire>
<wire>
<ID>1104 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-182,154,-182</points>
<connection>
<GID>836</GID>
<name>OUT_4</name></connection>
<connection>
<GID>875</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>930 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-138,105.5,-138</points>
<connection>
<GID>861</GID>
<name>OUT_3</name></connection>
<connection>
<GID>863</GID>
<name>IN_3</name></connection>
<intersection>98.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>98.5,-138,98.5,-124.5</points>
<connection>
<GID>951</GID>
<name>IN_0</name></connection>
<intersection>-138 1</intersection></vsegment></shape></wire>
<wire>
<ID>1107 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-180,154,-180</points>
<connection>
<GID>836</GID>
<name>OUT_6</name></connection>
<connection>
<GID>875</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1108 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-179,154,-179</points>
<connection>
<GID>836</GID>
<name>OUT_7</name></connection>
<connection>
<GID>875</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>891 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-96,105,-96</points>
<connection>
<GID>857</GID>
<name>OUT_12</name></connection>
<connection>
<GID>859</GID>
<name>IN_12</name></connection>
<intersection>80 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>80,-96,80,-91</points>
<connection>
<GID>942</GID>
<name>IN_0</name></connection>
<intersection>-96 1</intersection></vsegment></shape></wire>
<wire>
<ID>1098 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-178,154,-178</points>
<connection>
<GID>836</GID>
<name>OUT_8</name></connection>
<connection>
<GID>874</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1095 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>153.5,-177,154,-177</points>
<connection>
<GID>836</GID>
<name>OUT_9</name></connection>
<connection>
<GID>874</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>781 782 783 784 785 786 787 788 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-22,77,12</points>
<connection>
<GID>837</GID>
<name>OUT</name></connection>
<intersection>-22 2</intersection>
<intersection>12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,12,86,12</points>
<connection>
<GID>843</GID>
<name>OUT</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-22,83.5,-22</points>
<connection>
<GID>849</GID>
<name>OUT</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>1122 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-177,164.5,-177</points>
<connection>
<GID>876</GID>
<name>IN_1</name></connection>
<connection>
<GID>878</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>755 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-91.5,107,-89.5</points>
<connection>
<GID>984</GID>
<name>IN_0</name></connection>
<connection>
<GID>859</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1137 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-174,179,-174</points>
<connection>
<GID>877</GID>
<name>IN_4</name></connection>
<connection>
<GID>879</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>988 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,13.5,40,14</points>
<connection>
<GID>838</GID>
<name>OUT_0</name></connection>
<intersection>13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,13.5,42,13.5</points>
<connection>
<GID>869</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>789 790 791 792 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-29.5,79,6</points>
<intersection>-29.5 1</intersection>
<intersection>6 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-29.5,83.5,-29.5</points>
<connection>
<GID>851</GID>
<name>OUT</name></connection>
<intersection>77 4</intersection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79,6,86,6</points>
<connection>
<GID>841</GID>
<name>OUT</name></connection>
<intersection>79 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>77,-29.5,77,-28</points>
<connection>
<GID>839</GID>
<name>OUT</name></connection>
<intersection>-29.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1125 1126 1127 1128 1129 1130 1131 1132 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>158,-182.5,175,-182.5</points>
<connection>
<GID>875</GID>
<name>OUT</name></connection>
<intersection>175 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>175,-182.5,175,-174.5</points>
<connection>
<GID>879</GID>
<name>OUT</name></connection>
<intersection>-182.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1164 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-144,69.5,-144</points>
<connection>
<GID>897</GID>
<name>IN_0</name></connection>
<intersection>69.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>69.5,-144,69.5,-143</points>
<connection>
<GID>861</GID>
<name>clear</name></connection>
<intersection>-144 1</intersection></vsegment></shape></wire>
<wire>
<ID>801 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-26.5,105.5,-9.5</points>
<connection>
<GID>847</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>845</GID>
<name>ENABLE_0</name></connection>
<intersection>-9.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>105.5,-9.5,107,-9.5</points>
<connection>
<GID>982</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>795 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-24.5,103.5,-24.5</points>
<connection>
<GID>849</GID>
<name>IN_1</name></connection>
<connection>
<GID>845</GID>
<name>IN_1</name></connection>
<intersection>97.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>97.5,-24.5,97.5,-7.5</points>
<connection>
<GID>906</GID>
<name>IN_0</name></connection>
<intersection>-24.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>799 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-23.5,103.5,-23.5</points>
<connection>
<GID>849</GID>
<name>IN_2</name></connection>
<connection>
<GID>845</GID>
<name>IN_2</name></connection>
<intersection>96.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>96.5,-23.5,96.5,-15.5</points>
<connection>
<GID>907</GID>
<name>IN_0</name></connection>
<intersection>-23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1156 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-99,63,-99</points>
<connection>
<GID>857</GID>
<name>IN_9</name></connection>
<connection>
<GID>886</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>793 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-22.5,103.5,-22.5</points>
<connection>
<GID>849</GID>
<name>IN_3</name></connection>
<connection>
<GID>845</GID>
<name>IN_3</name></connection>
<intersection>95.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>95.5,-22.5,95.5,-7.5</points>
<connection>
<GID>908</GID>
<name>IN_0</name></connection>
<intersection>-22.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>798 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-21.5,103.5,-21.5</points>
<connection>
<GID>849</GID>
<name>IN_4</name></connection>
<connection>
<GID>845</GID>
<name>IN_4</name></connection>
<intersection>94.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>94.5,-21.5,94.5,-15.5</points>
<connection>
<GID>909</GID>
<name>IN_0</name></connection>
<intersection>-21.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>797 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-20.5,103.5,-20.5</points>
<connection>
<GID>849</GID>
<name>IN_5</name></connection>
<connection>
<GID>845</GID>
<name>IN_5</name></connection>
<intersection>93.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>93.5,-20.5,93.5,-7.5</points>
<connection>
<GID>910</GID>
<name>IN_0</name></connection>
<intersection>-20.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>794 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-19.5,103.5,-19.5</points>
<connection>
<GID>849</GID>
<name>IN_6</name></connection>
<connection>
<GID>845</GID>
<name>IN_6</name></connection>
<intersection>92.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>92.5,-19.5,92.5,-15.5</points>
<connection>
<GID>911</GID>
<name>IN_0</name></connection>
<intersection>-19.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1133 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-178,179,-178</points>
<connection>
<GID>877</GID>
<name>IN_0</name></connection>
<connection>
<GID>879</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>800 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-18.5,103.5,-18.5</points>
<connection>
<GID>849</GID>
<name>IN_7</name></connection>
<connection>
<GID>845</GID>
<name>IN_7</name></connection>
<intersection>91.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>91.5,-18.5,91.5,-7.5</points>
<connection>
<GID>912</GID>
<name>IN_0</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>839 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-26.5,107.5,-25.5</points>
<connection>
<GID>845</GID>
<name>OUT_0</name></connection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-26.5,110.5,-26.5</points>
<connection>
<GID>855</GID>
<name>IN_4</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>841 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-24.5,108.5,-23.5</points>
<intersection>-24.5 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-23.5,108.5,-23.5</points>
<connection>
<GID>845</GID>
<name>OUT_2</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,-24.5,110.5,-24.5</points>
<connection>
<GID>855</GID>
<name>IN_6</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1147 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-104,63,-104</points>
<connection>
<GID>857</GID>
<name>IN_4</name></connection>
<connection>
<GID>858</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>842 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,-23.5,109,-22.5</points>
<intersection>-23.5 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-22.5,109,-22.5</points>
<connection>
<GID>845</GID>
<name>OUT_3</name></connection>
<intersection>109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109,-23.5,110.5,-23.5</points>
<connection>
<GID>855</GID>
<name>IN_7</name></connection>
<intersection>109 0</intersection></hsegment></shape></wire>
<wire>
<ID>1178 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-91,68,-88.5</points>
<connection>
<GID>857</GID>
<name>count_enable</name></connection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-88.5,68,-88.5</points>
<connection>
<GID>952</GID>
<name>IN_0</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>843 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-22.5,109.5,-21.5</points>
<intersection>-22.5 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-21.5,109.5,-21.5</points>
<connection>
<GID>845</GID>
<name>OUT_4</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,-22.5,110.5,-22.5</points>
<connection>
<GID>855</GID>
<name>IN_8</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>844 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-21.5,110,-21</points>
<intersection>-21.5 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-21,110,-21</points>
<intersection>107.5 3</intersection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-21.5,110.5,-21.5</points>
<connection>
<GID>855</GID>
<name>IN_9</name></connection>
<intersection>110 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>107.5,-21,107.5,-20.5</points>
<connection>
<GID>845</GID>
<name>OUT_5</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>846 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-19.5,110,-19</points>
<intersection>-19.5 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-19,110,-19</points>
<intersection>107.5 3</intersection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-19.5,110.5,-19.5</points>
<connection>
<GID>855</GID>
<name>IN_11</name></connection>
<intersection>110 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>107.5,-19,107.5,-18.5</points>
<connection>
<GID>845</GID>
<name>OUT_7</name></connection>
<intersection>-19 1</intersection></vsegment></shape></wire>
<wire>
<ID>802 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-31,103.5,-31</points>
<connection>
<GID>851</GID>
<name>IN_0</name></connection>
<connection>
<GID>847</GID>
<name>IN_0</name></connection>
<intersection>102.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>102.5,-31,102.5,-15.5</points>
<connection>
<GID>901</GID>
<name>IN_0</name></connection>
<intersection>-31 1</intersection></vsegment></shape></wire>
<wire>
<ID>805 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-30,103.5,-30</points>
<connection>
<GID>851</GID>
<name>IN_1</name></connection>
<connection>
<GID>847</GID>
<name>IN_1</name></connection>
<intersection>101.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>101.5,-30,101.5,-7.5</points>
<connection>
<GID>902</GID>
<name>IN_0</name></connection>
<intersection>-30 1</intersection></vsegment></shape></wire>
<wire>
<ID>1138 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-172,179,-172</points>
<connection>
<GID>877</GID>
<name>IN_6</name></connection>
<connection>
<GID>879</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>803 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-29,103.5,-29</points>
<connection>
<GID>851</GID>
<name>IN_2</name></connection>
<connection>
<GID>847</GID>
<name>IN_2</name></connection>
<intersection>100.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>100.5,-29,100.5,-15.5</points>
<connection>
<GID>903</GID>
<name>IN_0</name></connection>
<intersection>-29 1</intersection></vsegment></shape></wire>
<wire>
<ID>804 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-28,103.5,-28</points>
<connection>
<GID>851</GID>
<name>IN_3</name></connection>
<connection>
<GID>847</GID>
<name>IN_3</name></connection>
<intersection>99.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>99.5,-28,99.5,-7.5</points>
<connection>
<GID>904</GID>
<name>IN_0</name></connection>
<intersection>-28 1</intersection></vsegment></shape></wire>
<wire>
<ID>836 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>107.5,-29.5,110.5,-29.5</points>
<connection>
<GID>855</GID>
<name>IN_1</name></connection>
<intersection>107.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>107.5,-30,107.5,-29.5</points>
<connection>
<GID>847</GID>
<name>OUT_1</name></connection>
<intersection>-29.5 0</intersection></vsegment></shape></wire>
<wire>
<ID>838 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>107.5,-27.5,110.5,-27.5</points>
<connection>
<GID>855</GID>
<name>IN_3</name></connection>
<intersection>107.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>107.5,-28,107.5,-27.5</points>
<connection>
<GID>847</GID>
<name>OUT_3</name></connection>
<intersection>-27.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>822 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-49.5,106,-40.5</points>
<connection>
<GID>854</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>853</GID>
<name>ENABLE_0</name></connection>
<intersection>-40.5 31</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>105,-40.5,106,-40.5</points>
<connection>
<GID>961</GID>
<name>IN_0</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>1150 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-98,63,-98</points>
<connection>
<GID>857</GID>
<name>IN_10</name></connection>
<connection>
<GID>887</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>978 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-166.5,111,-166.5</points>
<connection>
<GID>866</GID>
<name>OUT_1</name></connection>
<connection>
<GID>865</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1155 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-97,63,-97</points>
<connection>
<GID>857</GID>
<name>IN_11</name></connection>
<connection>
<GID>888</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1151 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-96,63,-96</points>
<connection>
<GID>857</GID>
<name>IN_12</name></connection>
<connection>
<GID>889</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>947 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-130,111,-130</points>
<connection>
<GID>863</GID>
<name>OUT_11</name></connection>
<connection>
<GID>862</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1154 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-95,63,-95</points>
<connection>
<GID>857</GID>
<name>IN_13</name></connection>
<connection>
<GID>890</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>973 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-160.5,111,-160.5</points>
<connection>
<GID>866</GID>
<name>OUT_7</name></connection>
<connection>
<GID>865</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1152 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-94,63,-94</points>
<connection>
<GID>857</GID>
<name>IN_14</name></connection>
<connection>
<GID>891</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1153 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-93,63,-93</points>
<connection>
<GID>857</GID>
<name>IN_15</name></connection>
<connection>
<GID>892</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1158 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-103,63,-103</points>
<connection>
<GID>857</GID>
<name>IN_5</name></connection>
<connection>
<GID>860</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1148 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-102,63,-102</points>
<connection>
<GID>857</GID>
<name>IN_6</name></connection>
<connection>
<GID>883</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>952 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-139,111,-139</points>
<connection>
<GID>863</GID>
<name>OUT_2</name></connection>
<connection>
<GID>862</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1157 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-101,63,-101</points>
<connection>
<GID>857</GID>
<name>IN_7</name></connection>
<connection>
<GID>884</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>986 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-167.5,111,-167.5</points>
<connection>
<GID>866</GID>
<name>OUT_0</name></connection>
<connection>
<GID>865</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1163 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>67,-112,69,-112</points>
<connection>
<GID>896</GID>
<name>IN_0</name></connection>
<intersection>69 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>69,-112,69,-110</points>
<connection>
<GID>857</GID>
<name>clear</name></connection>
<intersection>-112 1</intersection></vsegment></shape></wire>
<wire>
<ID>1177 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-91,67,-90.5</points>
<connection>
<GID>857</GID>
<name>load</name></connection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-90.5,67,-90.5</points>
<connection>
<GID>975</GID>
<name>IN_0</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>899 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-108,105,-108</points>
<connection>
<GID>857</GID>
<name>OUT_0</name></connection>
<connection>
<GID>859</GID>
<name>IN_0</name></connection>
<intersection>104 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>104,-108,104,-91</points>
<connection>
<GID>929</GID>
<name>IN_0</name></connection>
<intersection>-108 1</intersection></vsegment></shape></wire>
<wire>
<ID>903 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-107,105,-107</points>
<connection>
<GID>857</GID>
<name>OUT_1</name></connection>
<connection>
<GID>859</GID>
<name>IN_1</name></connection>
<intersection>102 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>102,-107,102,-91</points>
<connection>
<GID>930</GID>
<name>IN_0</name></connection>
<intersection>-107 1</intersection></vsegment></shape></wire>
<wire>
<ID>896 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-98,105,-98</points>
<connection>
<GID>857</GID>
<name>OUT_10</name></connection>
<connection>
<GID>859</GID>
<name>IN_10</name></connection>
<intersection>84 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>84,-98,84,-91</points>
<connection>
<GID>939</GID>
<name>IN_0</name></connection>
<intersection>-98 1</intersection></vsegment></shape></wire>
<wire>
<ID>902 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-97,105,-97</points>
<connection>
<GID>857</GID>
<name>OUT_11</name></connection>
<connection>
<GID>859</GID>
<name>IN_11</name></connection>
<intersection>82 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>82,-97,82,-91</points>
<connection>
<GID>941</GID>
<name>IN_0</name></connection>
<intersection>-97 1</intersection></vsegment></shape></wire>
<wire>
<ID>892 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-95,105,-95</points>
<connection>
<GID>857</GID>
<name>OUT_13</name></connection>
<connection>
<GID>859</GID>
<name>IN_13</name></connection>
<intersection>78 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>78,-95,78,-91</points>
<connection>
<GID>943</GID>
<name>IN_0</name></connection>
<intersection>-95 1</intersection></vsegment></shape></wire>
<wire>
<ID>905 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-94,105,-94</points>
<connection>
<GID>857</GID>
<name>OUT_14</name></connection>
<connection>
<GID>859</GID>
<name>IN_14</name></connection>
<intersection>76 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>76,-94,76,-91</points>
<connection>
<GID>944</GID>
<name>IN_0</name></connection>
<intersection>-94 1</intersection></vsegment></shape></wire>
<wire>
<ID>906 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-93,105,-93</points>
<connection>
<GID>857</GID>
<name>OUT_15</name></connection>
<connection>
<GID>859</GID>
<name>IN_15</name></connection>
<intersection>74 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>74,-93,74,-91</points>
<connection>
<GID>945</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>897 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-106,105,-106</points>
<connection>
<GID>857</GID>
<name>OUT_2</name></connection>
<connection>
<GID>859</GID>
<name>IN_2</name></connection>
<intersection>100 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>100,-106,100,-91</points>
<connection>
<GID>931</GID>
<name>IN_0</name></connection>
<intersection>-106 1</intersection></vsegment></shape></wire>
<wire>
<ID>898 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-105,105,-105</points>
<connection>
<GID>857</GID>
<name>OUT_3</name></connection>
<connection>
<GID>859</GID>
<name>IN_3</name></connection>
<intersection>98 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>98,-105,98,-91</points>
<connection>
<GID>932</GID>
<name>IN_0</name></connection>
<intersection>-105 1</intersection></vsegment></shape></wire>
<wire>
<ID>1049 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-156.5,63.5,-156.5</points>
<connection>
<GID>871</GID>
<name>IN_11</name></connection>
<connection>
<GID>864</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>900 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-104,105,-104</points>
<connection>
<GID>857</GID>
<name>OUT_4</name></connection>
<connection>
<GID>859</GID>
<name>IN_4</name></connection>
<intersection>96 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>96,-104,96,-91</points>
<connection>
<GID>933</GID>
<name>IN_0</name></connection>
<intersection>-104 1</intersection></vsegment></shape></wire>
<wire>
<ID>894 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-103,105,-103</points>
<connection>
<GID>857</GID>
<name>OUT_5</name></connection>
<connection>
<GID>859</GID>
<name>IN_5</name></connection>
<intersection>94 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>94,-103,94,-91</points>
<connection>
<GID>934</GID>
<name>IN_0</name></connection>
<intersection>-103 1</intersection></vsegment></shape></wire>
<wire>
<ID>901 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-102,105,-102</points>
<connection>
<GID>857</GID>
<name>OUT_6</name></connection>
<connection>
<GID>859</GID>
<name>IN_6</name></connection>
<intersection>92 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>92,-102,92,-91</points>
<connection>
<GID>935</GID>
<name>IN_0</name></connection>
<intersection>-102 1</intersection></vsegment></shape></wire>
<wire>
<ID>904 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-101,105,-101</points>
<connection>
<GID>857</GID>
<name>OUT_7</name></connection>
<connection>
<GID>859</GID>
<name>IN_7</name></connection>
<intersection>90 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>90,-101,90,-91</points>
<connection>
<GID>936</GID>
<name>IN_0</name></connection>
<intersection>-101 1</intersection></vsegment></shape></wire>
<wire>
<ID>895 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-100,105,-100</points>
<connection>
<GID>857</GID>
<name>OUT_8</name></connection>
<connection>
<GID>859</GID>
<name>IN_8</name></connection>
<intersection>88 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>88,-100,88,-91</points>
<connection>
<GID>937</GID>
<name>IN_0</name></connection>
<intersection>-100 1</intersection></vsegment></shape></wire>
<wire>
<ID>1036 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-131,63.5,-131</points>
<connection>
<GID>870</GID>
<name>IN_10</name></connection>
<connection>
<GID>861</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1042 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-129,63.5,-129</points>
<connection>
<GID>870</GID>
<name>IN_12</name></connection>
<connection>
<GID>861</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1044 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-127,63.5,-127</points>
<connection>
<GID>870</GID>
<name>IN_14</name></connection>
<connection>
<GID>861</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1037 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-138,63.5,-138</points>
<connection>
<GID>870</GID>
<name>IN_3</name></connection>
<connection>
<GID>861</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1038 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-137,63.5,-137</points>
<connection>
<GID>870</GID>
<name>IN_4</name></connection>
<connection>
<GID>861</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1039 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-136,63.5,-136</points>
<connection>
<GID>870</GID>
<name>IN_5</name></connection>
<connection>
<GID>861</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1031 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-135,63.5,-135</points>
<connection>
<GID>870</GID>
<name>IN_6</name></connection>
<connection>
<GID>861</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1030 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-134,63.5,-134</points>
<connection>
<GID>870</GID>
<name>IN_7</name></connection>
<connection>
<GID>861</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1182 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-124,69.5,-118.5</points>
<connection>
<GID>861</GID>
<name>count_up</name></connection>
<intersection>-118.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-118.5,69.5,-118.5</points>
<connection>
<GID>958</GID>
<name>IN_0</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>931 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-141,105.5,-141</points>
<connection>
<GID>861</GID>
<name>OUT_0</name></connection>
<connection>
<GID>863</GID>
<name>IN_0</name></connection>
<intersection>104.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>104.5,-141,104.5,-124.5</points>
<connection>
<GID>947</GID>
<name>IN_0</name></connection>
<intersection>-141 1</intersection></vsegment></shape></wire>
<wire>
<ID>935 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-140,105.5,-140</points>
<connection>
<GID>861</GID>
<name>OUT_1</name></connection>
<connection>
<GID>863</GID>
<name>IN_1</name></connection>
<intersection>102.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>102.5,-140,102.5,-124.5</points>
<connection>
<GID>948</GID>
<name>IN_0</name></connection>
<intersection>-140 1</intersection></vsegment></shape></wire>
<wire>
<ID>928 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-131,105.5,-131</points>
<connection>
<GID>861</GID>
<name>OUT_10</name></connection>
<connection>
<GID>863</GID>
<name>IN_10</name></connection>
<intersection>84.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>84.5,-131,84.5,-124.5</points>
<connection>
<GID>962</GID>
<name>IN_0</name></connection>
<intersection>-131 1</intersection></vsegment></shape></wire>
<wire>
<ID>934 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-130,105.5,-130</points>
<connection>
<GID>861</GID>
<name>OUT_11</name></connection>
<connection>
<GID>863</GID>
<name>IN_11</name></connection>
<intersection>82.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>82.5,-130,82.5,-124.5</points>
<connection>
<GID>963</GID>
<name>IN_0</name></connection>
<intersection>-130 1</intersection></vsegment></shape></wire>
<wire>
<ID>923 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-129,105.5,-129</points>
<connection>
<GID>861</GID>
<name>OUT_12</name></connection>
<connection>
<GID>863</GID>
<name>IN_12</name></connection>
<intersection>80.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>80.5,-129,80.5,-124.5</points>
<connection>
<GID>964</GID>
<name>IN_0</name></connection>
<intersection>-129 1</intersection></vsegment></shape></wire>
<wire>
<ID>937 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-127,105.5,-127</points>
<connection>
<GID>861</GID>
<name>OUT_14</name></connection>
<connection>
<GID>863</GID>
<name>IN_14</name></connection>
<intersection>76.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>76.5,-127,76.5,-124.5</points>
<connection>
<GID>967</GID>
<name>IN_0</name></connection>
<intersection>-127 1</intersection></vsegment></shape></wire>
<wire>
<ID>938 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-126,105.5,-126</points>
<connection>
<GID>861</GID>
<name>OUT_15</name></connection>
<connection>
<GID>863</GID>
<name>IN_15</name></connection>
<intersection>74.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>74.5,-126,74.5,-124.5</points>
<connection>
<GID>968</GID>
<name>IN_0</name></connection>
<intersection>-126 1</intersection></vsegment></shape></wire>
<wire>
<ID>929 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-139,105.5,-139</points>
<connection>
<GID>861</GID>
<name>OUT_2</name></connection>
<connection>
<GID>863</GID>
<name>IN_2</name></connection>
<intersection>100.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>100.5,-139,100.5,-124.5</points>
<connection>
<GID>950</GID>
<name>IN_0</name></connection>
<intersection>-139 1</intersection></vsegment></shape></wire>
<wire>
<ID>926 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-136,105.5,-136</points>
<connection>
<GID>861</GID>
<name>OUT_5</name></connection>
<connection>
<GID>863</GID>
<name>IN_5</name></connection>
<intersection>94.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>94.5,-136,94.5,-124.5</points>
<connection>
<GID>954</GID>
<name>IN_0</name></connection>
<intersection>-136 1</intersection></vsegment></shape></wire>
<wire>
<ID>933 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-135,105.5,-135</points>
<connection>
<GID>861</GID>
<name>OUT_6</name></connection>
<connection>
<GID>863</GID>
<name>IN_6</name></connection>
<intersection>92.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>92.5,-135,92.5,-124.5</points>
<connection>
<GID>956</GID>
<name>IN_0</name></connection>
<intersection>-135 1</intersection></vsegment></shape></wire>
<wire>
<ID>936 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-134,105.5,-134</points>
<connection>
<GID>861</GID>
<name>OUT_7</name></connection>
<connection>
<GID>863</GID>
<name>IN_7</name></connection>
<intersection>90.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>90.5,-134,90.5,-124.5</points>
<connection>
<GID>957</GID>
<name>IN_0</name></connection>
<intersection>-134 1</intersection></vsegment></shape></wire>
<wire>
<ID>927 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-133,105.5,-133</points>
<connection>
<GID>861</GID>
<name>OUT_8</name></connection>
<connection>
<GID>863</GID>
<name>IN_8</name></connection>
<intersection>88.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>88.5,-133,88.5,-124.5</points>
<connection>
<GID>959</GID>
<name>IN_0</name></connection>
<intersection>-133 1</intersection></vsegment></shape></wire>
<wire>
<ID>954 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-141,111,-141</points>
<connection>
<GID>863</GID>
<name>OUT_0</name></connection>
<connection>
<GID>862</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1123 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-171,164.5,-171</points>
<connection>
<GID>876</GID>
<name>IN_7</name></connection>
<connection>
<GID>878</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>946 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-140,111,-140</points>
<connection>
<GID>863</GID>
<name>OUT_1</name></connection>
<connection>
<GID>862</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>945 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-131,111,-131</points>
<connection>
<GID>863</GID>
<name>OUT_10</name></connection>
<connection>
<GID>862</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>948 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-129,111,-129</points>
<connection>
<GID>863</GID>
<name>OUT_12</name></connection>
<connection>
<GID>862</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>943 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-128,111,-128</points>
<connection>
<GID>863</GID>
<name>OUT_13</name></connection>
<connection>
<GID>862</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>951 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-127,111,-127</points>
<connection>
<GID>863</GID>
<name>OUT_14</name></connection>
<connection>
<GID>862</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>950 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-126,111,-126</points>
<connection>
<GID>863</GID>
<name>OUT_15</name></connection>
<connection>
<GID>862</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>944 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-138,111,-138</points>
<connection>
<GID>863</GID>
<name>OUT_3</name></connection>
<connection>
<GID>862</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>940 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-137,111,-137</points>
<connection>
<GID>863</GID>
<name>OUT_4</name></connection>
<connection>
<GID>862</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>939 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-136,111,-136</points>
<connection>
<GID>863</GID>
<name>OUT_5</name></connection>
<connection>
<GID>862</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>942 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-135,111,-135</points>
<connection>
<GID>863</GID>
<name>OUT_6</name></connection>
<connection>
<GID>862</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1120 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-173,164.5,-173</points>
<connection>
<GID>876</GID>
<name>IN_5</name></connection>
<connection>
<GID>878</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>941 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-134,111,-134</points>
<connection>
<GID>863</GID>
<name>OUT_7</name></connection>
<connection>
<GID>862</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>953 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-133,111,-133</points>
<connection>
<GID>863</GID>
<name>OUT_8</name></connection>
<connection>
<GID>862</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>949 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-132,111,-132</points>
<connection>
<GID>863</GID>
<name>OUT_9</name></connection>
<connection>
<GID>862</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>756 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-124.5,107.5,-121.5</points>
<connection>
<GID>985</GID>
<name>IN_0</name></connection>
<connection>
<GID>863</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1045 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-167.5,63.5,-167.5</points>
<connection>
<GID>871</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>864</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1055 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-155.5,63.5,-155.5</points>
<connection>
<GID>871</GID>
<name>IN_12</name></connection>
<connection>
<GID>864</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1050 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-154.5,63.5,-154.5</points>
<connection>
<GID>871</GID>
<name>IN_13</name></connection>
<connection>
<GID>864</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1060 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-152.5,63.5,-152.5</points>
<connection>
<GID>871</GID>
<name>IN_15</name></connection>
<connection>
<GID>864</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1047 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-165.5,63.5,-165.5</points>
<connection>
<GID>871</GID>
<name>IN_2</name></connection>
<connection>
<GID>864</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1046 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-163.5,63.5,-163.5</points>
<connection>
<GID>871</GID>
<name>IN_4</name></connection>
<connection>
<GID>864</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1052 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-161.5,63.5,-161.5</points>
<connection>
<GID>871</GID>
<name>IN_6</name></connection>
<connection>
<GID>864</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1054 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-160.5,63.5,-160.5</points>
<connection>
<GID>871</GID>
<name>IN_7</name></connection>
<connection>
<GID>864</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1053 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-159.5,63.5,-159.5</points>
<connection>
<GID>871</GID>
<name>IN_8</name></connection>
<connection>
<GID>864</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1058 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-158.5,63.5,-158.5</points>
<connection>
<GID>871</GID>
<name>IN_9</name></connection>
<connection>
<GID>864</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1185 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-150.5,69.5,-146</points>
<connection>
<GID>864</GID>
<name>count_up</name></connection>
<intersection>-146 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-146,69.5,-146</points>
<connection>
<GID>979</GID>
<name>IN_0</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1183 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-150.5,67.5,-150</points>
<connection>
<GID>864</GID>
<name>load</name></connection>
<intersection>-150 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-150,67.5,-150</points>
<connection>
<GID>978</GID>
<name>IN_0</name></connection>
<intersection>67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>963 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-167.5,104,-167.5</points>
<connection>
<GID>864</GID>
<name>OUT_0</name></connection>
<connection>
<GID>866</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>960 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-157.5,104,-157.5</points>
<connection>
<GID>864</GID>
<name>OUT_10</name></connection>
<connection>
<GID>866</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>966 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-156.5,104,-156.5</points>
<connection>
<GID>864</GID>
<name>OUT_11</name></connection>
<connection>
<GID>866</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>956 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-154.5,104,-154.5</points>
<connection>
<GID>864</GID>
<name>OUT_13</name></connection>
<connection>
<GID>866</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>969 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-153.5,104,-153.5</points>
<connection>
<GID>864</GID>
<name>OUT_14</name></connection>
<connection>
<GID>866</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>970 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-152.5,104,-152.5</points>
<connection>
<GID>864</GID>
<name>OUT_15</name></connection>
<connection>
<GID>866</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>961 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-165.5,104,-165.5</points>
<connection>
<GID>864</GID>
<name>OUT_2</name></connection>
<connection>
<GID>866</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>962 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-164.5,104,-164.5</points>
<connection>
<GID>864</GID>
<name>OUT_3</name></connection>
<connection>
<GID>866</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>964 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-163.5,104,-163.5</points>
<connection>
<GID>864</GID>
<name>OUT_4</name></connection>
<connection>
<GID>866</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>958 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-162.5,104,-162.5</points>
<connection>
<GID>864</GID>
<name>OUT_5</name></connection>
<connection>
<GID>866</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>965 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-161.5,104,-161.5</points>
<connection>
<GID>864</GID>
<name>OUT_6</name></connection>
<connection>
<GID>866</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>968 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-160.5,104,-160.5</points>
<connection>
<GID>864</GID>
<name>OUT_7</name></connection>
<connection>
<GID>866</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>959 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-159.5,104,-159.5</points>
<connection>
<GID>864</GID>
<name>OUT_8</name></connection>
<connection>
<GID>866</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1136 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-175,179,-175</points>
<connection>
<GID>877</GID>
<name>IN_3</name></connection>
<connection>
<GID>879</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>957 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-158.5,104,-158.5</points>
<connection>
<GID>864</GID>
<name>OUT_9</name></connection>
<connection>
<GID>866</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>977 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-157.5,111,-157.5</points>
<connection>
<GID>866</GID>
<name>OUT_10</name></connection>
<connection>
<GID>865</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>979 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-156.5,111,-156.5</points>
<connection>
<GID>866</GID>
<name>OUT_11</name></connection>
<connection>
<GID>865</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>980 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-155.5,111,-155.5</points>
<connection>
<GID>866</GID>
<name>OUT_12</name></connection>
<connection>
<GID>865</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>975 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-154.5,111,-154.5</points>
<connection>
<GID>866</GID>
<name>OUT_13</name></connection>
<connection>
<GID>865</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>983 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-153.5,111,-153.5</points>
<connection>
<GID>866</GID>
<name>OUT_14</name></connection>
<connection>
<GID>865</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>982 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-152.5,111,-152.5</points>
<connection>
<GID>866</GID>
<name>OUT_15</name></connection>
<connection>
<GID>865</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>984 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-165.5,111,-165.5</points>
<connection>
<GID>866</GID>
<name>OUT_2</name></connection>
<connection>
<GID>865</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>976 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-164.5,111,-164.5</points>
<connection>
<GID>866</GID>
<name>OUT_3</name></connection>
<connection>
<GID>865</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1121 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-174,164.5,-174</points>
<connection>
<GID>876</GID>
<name>IN_4</name></connection>
<connection>
<GID>878</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>972 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-163.5,111,-163.5</points>
<connection>
<GID>866</GID>
<name>OUT_4</name></connection>
<connection>
<GID>865</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>971 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-162.5,111,-162.5</points>
<connection>
<GID>866</GID>
<name>OUT_5</name></connection>
<connection>
<GID>865</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>974 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-161.5,111,-161.5</points>
<connection>
<GID>866</GID>
<name>OUT_6</name></connection>
<connection>
<GID>865</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>985 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-159.5,111,-159.5</points>
<connection>
<GID>866</GID>
<name>OUT_8</name></connection>
<connection>
<GID>865</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1119 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-178,164.5,-178</points>
<connection>
<GID>876</GID>
<name>IN_0</name></connection>
<connection>
<GID>878</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1124 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-175,164.5,-175</points>
<connection>
<GID>876</GID>
<name>IN_3</name></connection>
<connection>
<GID>878</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>1134 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-177,179,-177</points>
<connection>
<GID>877</GID>
<name>IN_1</name></connection>
<connection>
<GID>879</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1135 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-176,179,-176</points>
<connection>
<GID>877</GID>
<name>IN_2</name></connection>
<connection>
<GID>879</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1140 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-171,179,-171</points>
<connection>
<GID>877</GID>
<name>IN_7</name></connection>
<connection>
<GID>879</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>1191 </ID>
<shape>
<hsegment>
<ID>4</ID>
<points>42,0,45,0</points>
<connection>
<GID>994</GID>
<name>IN_0</name></connection>
<connection>
<GID>990</GID>
<name>OUT_0</name></connection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-72.9287,1232.88,1323.07,549.883</PageViewport></page 3></circuit>