
<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-32.95,39.6893,61.95,-63.2229</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>14.5,-13</position>
<gparam>LABEL_TEXT Go to https://cedar.to/vjyQw7 to download the latest version!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>14.5,-9.5</position>
<gparam>LABEL_TEXT Error: This file was made with a newer version of Cedar Logic!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate></page 0>
</circuit>
<throw_away></throw_away>

	<version>2.3 | 2018-03- 4 22:33:02</version><circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-18.896,9.8258,156.842,-76.1548</PageViewport>
<gate>
<ID>70</ID>
<type>BW_8X1_BUS_END</type>
<position>92,-34</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>166 </input>
<input>
<ID>IN_2</ID>167 </input>
<input>
<ID>IN_3</ID>164 </input>
<input>
<ID>IN_4</ID>169 </input>
<input>
<ID>IN_5</ID>168 </input>
<input>
<ID>IN_6</ID>170 </input>
<input>
<ID>IN_7</ID>171 </input>
<input>
<ID>OUT</ID>81 82 83 84 85 86 87 88 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>6</ID>
<type>BI_ROM_12x16</type>
<position>25,-17</position>
<input>
<ID>ADDRESS_0</ID>130 </input>
<input>
<ID>ADDRESS_1</ID>125 </input>
<input>
<ID>ADDRESS_2</ID>131 </input>
<input>
<ID>ADDRESS_3</ID>124 </input>
<input>
<ID>ADDRESS_4</ID>127 </input>
<input>
<ID>ADDRESS_5</ID>126 </input>
<input>
<ID>ADDRESS_6</ID>129 </input>
<input>
<ID>ADDRESS_7</ID>128 </input>
<output>
<ID>DATA_OUT_0</ID>28 </output>
<output>
<ID>DATA_OUT_1</ID>27 </output>
<output>
<ID>DATA_OUT_10</ID>112 </output>
<output>
<ID>DATA_OUT_11</ID>113 </output>
<output>
<ID>DATA_OUT_12</ID>114 </output>
<output>
<ID>DATA_OUT_13</ID>115 </output>
<output>
<ID>DATA_OUT_14</ID>185 </output>
<output>
<ID>DATA_OUT_15</ID>186 </output>
<output>
<ID>DATA_OUT_2</ID>26 </output>
<output>
<ID>DATA_OUT_3</ID>31 </output>
<output>
<ID>DATA_OUT_4</ID>29 </output>
<output>
<ID>DATA_OUT_5</ID>30 </output>
<output>
<ID>DATA_OUT_6</ID>32 </output>
<output>
<ID>DATA_OUT_7</ID>25 </output>
<output>
<ID>DATA_OUT_8</ID>110 </output>
<output>
<ID>DATA_OUT_9</ID>111 </output>
<input>
<ID>ENABLE_0</ID>183 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:0 4352</lparam>
<lparam>Address:2 513</lparam>
<lparam>Address:3 5632</lparam>
<lparam>Address:5 769</lparam></gate>
<gate>
<ID>86</ID>
<type>EE_VDD</type>
<position>35,-13.5</position>
<output>
<ID>OUT_0</ID>183 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>22</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>45.5,-34.5</position>
<input>
<ID>ENABLE_0</ID>180 </input>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>63 </input>
<input>
<ID>IN_3</ID>62 </input>
<input>
<ID>IN_4</ID>60 </input>
<input>
<ID>IN_5</ID>64 </input>
<input>
<ID>IN_6</ID>59 </input>
<input>
<ID>IN_7</ID>61 </input>
<output>
<ID>OUT_0</ID>67 </output>
<output>
<ID>OUT_1</ID>66 </output>
<output>
<ID>OUT_2</ID>72 </output>
<output>
<ID>OUT_3</ID>65 </output>
<output>
<ID>OUT_4</ID>68 </output>
<output>
<ID>OUT_5</ID>69 </output>
<output>
<ID>OUT_6</ID>71 </output>
<output>
<ID>OUT_7</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>9</ID>
<type>BW_8X1_BUS_END</type>
<position>29,-31</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>27 </input>
<input>
<ID>IN_2</ID>26 </input>
<input>
<ID>IN_3</ID>31 </input>
<input>
<ID>IN_4</ID>29 </input>
<input>
<ID>IN_5</ID>30 </input>
<input>
<ID>IN_6</ID>32 </input>
<input>
<ID>IN_7</ID>25 </input>
<input>
<ID>OUT</ID>49 50 51 52 53 54 55 56 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>84</ID>
<type>DA_FROM</type>
<position>59,-9.5</position>
<input>
<ID>IN_0</ID>182 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>20</ID>
<type>BW_8X1_BUS_END</type>
<position>41.5,-34.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>63 </input>
<input>
<ID>IN_3</ID>62 </input>
<input>
<ID>IN_4</ID>60 </input>
<input>
<ID>IN_5</ID>64 </input>
<input>
<ID>IN_6</ID>59 </input>
<input>
<ID>IN_7</ID>61 </input>
<input>
<ID>OUT</ID>49 50 51 52 53 54 55 56 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>47,-27</position>
<input>
<ID>IN_0</ID>180 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Pass_value</lparam></gate>
<gate>
<ID>18</ID>
<type>AE_RAM_8x8</type>
<position>56.5,-16.5</position>
<input>
<ID>ADDRESS_0</ID>41 </input>
<input>
<ID>ADDRESS_1</ID>46 </input>
<input>
<ID>ADDRESS_2</ID>47 </input>
<input>
<ID>ADDRESS_3</ID>45 </input>
<input>
<ID>ADDRESS_4</ID>48 </input>
<input>
<ID>ADDRESS_5</ID>42 </input>
<input>
<ID>ADDRESS_6</ID>43 </input>
<input>
<ID>ADDRESS_7</ID>44 </input>
<input>
<ID>DATA_IN_0</ID>73 </input>
<input>
<ID>DATA_IN_1</ID>77 </input>
<input>
<ID>DATA_IN_2</ID>78 </input>
<input>
<ID>DATA_IN_3</ID>74 </input>
<input>
<ID>DATA_IN_4</ID>79 </input>
<input>
<ID>DATA_IN_5</ID>80 </input>
<input>
<ID>DATA_IN_6</ID>75 </input>
<input>
<ID>DATA_IN_7</ID>76 </input>
<output>
<ID>DATA_OUT_0</ID>73 </output>
<output>
<ID>DATA_OUT_1</ID>77 </output>
<output>
<ID>DATA_OUT_2</ID>78 </output>
<output>
<ID>DATA_OUT_3</ID>74 </output>
<output>
<ID>DATA_OUT_4</ID>79 </output>
<output>
<ID>DATA_OUT_5</ID>80 </output>
<output>
<ID>DATA_OUT_6</ID>75 </output>
<output>
<ID>DATA_OUT_7</ID>76 </output>
<input>
<ID>ENABLE_0</ID>179 </input>
<input>
<ID>write_clock</ID>182 </input>
<input>
<ID>write_enable</ID>181 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:0 5</lparam>
<lparam>Address:1 2</lparam>
<lparam>Address:2 35</lparam></gate>
<gate>
<ID>19</ID>
<type>BW_8X1_BUS_END</type>
<position>48.5,-16.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>46 </input>
<input>
<ID>IN_2</ID>47 </input>
<input>
<ID>IN_3</ID>45 </input>
<input>
<ID>IN_4</ID>48 </input>
<input>
<ID>IN_5</ID>42 </input>
<input>
<ID>IN_6</ID>43 </input>
<input>
<ID>IN_7</ID>44 </input>
<input>
<ID>OUT</ID>49 50 51 52 53 54 55 56 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>59,-7</position>
<input>
<ID>IN_0</ID>181 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID write</lparam></gate>
<gate>
<ID>24</ID>
<type>BW_8X1_BUS_END</type>
<position>49.5,-34.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>66 </input>
<input>
<ID>IN_2</ID>72 </input>
<input>
<ID>IN_3</ID>65 </input>
<input>
<ID>IN_4</ID>68 </input>
<input>
<ID>IN_5</ID>69 </input>
<input>
<ID>IN_6</ID>71 </input>
<input>
<ID>IN_7</ID>70 </input>
<input>
<ID>OUT</ID>81 82 83 84 85 86 87 88 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>88</ID>
<type>DA_FROM</type>
<position>72.5,-12</position>
<input>
<ID>IN_0</ID>184 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C4</lparam></gate>
<gate>
<ID>25</ID>
<type>BW_8X1_BUS_END</type>
<position>56.5,-25.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>77 </input>
<input>
<ID>IN_2</ID>78 </input>
<input>
<ID>IN_3</ID>74 </input>
<input>
<ID>IN_4</ID>79 </input>
<input>
<ID>IN_5</ID>80 </input>
<input>
<ID>IN_6</ID>75 </input>
<input>
<ID>IN_7</ID>76 </input>
<input>
<ID>OUT</ID>81 82 83 84 85 86 87 88 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>89</ID>
<type>DE_TO</type>
<position>31,-43.5</position>
<input>
<ID>IN_0</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C6</lparam></gate>
<gate>
<ID>27</ID>
<type>BW_8X1_BUS_END</type>
<position>100.5,-34.5</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>99 </input>
<input>
<ID>IN_2</ID>100 </input>
<input>
<ID>IN_3</ID>101 </input>
<input>
<ID>IN_4</ID>102 </input>
<input>
<ID>IN_5</ID>103 </input>
<input>
<ID>IN_6</ID>13 </input>
<input>
<ID>IN_7</ID>14 </input>
<input>
<ID>OUT</ID>81 82 83 84 85 86 87 88 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>91</ID>
<type>DA_FROM</type>
<position>80,-25</position>
<input>
<ID>IN_0</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_REGISTER8</type>
<position>83,-19</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>91 </input>
<input>
<ID>IN_2</ID>94 </input>
<input>
<ID>IN_3</ID>92 </input>
<input>
<ID>IN_4</ID>97 </input>
<input>
<ID>IN_5</ID>96 </input>
<input>
<ID>IN_6</ID>11 </input>
<input>
<ID>IN_7</ID>12 </input>
<output>
<ID>OUT_0</ID>104 </output>
<output>
<ID>OUT_1</ID>105 </output>
<output>
<ID>OUT_2</ID>106 </output>
<output>
<ID>OUT_3</ID>107 </output>
<output>
<ID>OUT_4</ID>108 </output>
<output>
<ID>OUT_5</ID>109 </output>
<output>
<ID>OUT_6</ID>6 </output>
<output>
<ID>OUT_7</ID>7 </output>
<input>
<ID>clock</ID>187 </input>
<input>
<ID>load</ID>184 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 5</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>71.5,-22</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>76.5,-21</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>71.5,-20</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R2</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>76.5,-19</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R3</lparam></gate>
<gate>
<ID>37</ID>
<type>DA_FROM</type>
<position>71.5,-18</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R4</lparam></gate>
<gate>
<ID>101</ID>
<type>CC_PULSE</type>
<position>-17.5,-1</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>DA_FROM</type>
<position>76.5,-17</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R5</lparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>106,-38</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>43</ID>
<type>DE_TO</type>
<position>111,-37</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>106,-36</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_TO</type>
<position>111,-35</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>106,-34</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>110</ID>
<type>DE_TO</type>
<position>-12,-3.5</position>
<input>
<ID>IN_0</ID>195 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>111,-33</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>100.5,-22</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_TOGGLE</type>
<position>-17.5,-3.5</position>
<output>
<ID>OUT_0</ID>195 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>DE_TO</type>
<position>105.5,-21</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>50</ID>
<type>DE_TO</type>
<position>100.5,-20</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>51</ID>
<type>DE_TO</type>
<position>105.5,-19</position>
<input>
<ID>IN_0</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>52</ID>
<type>DE_TO</type>
<position>100.5,-18</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>53</ID>
<type>DE_TO</type>
<position>105.5,-17</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>55</ID>
<type>DE_TO</type>
<position>31,-55.5</position>
<input>
<ID>IN_0</ID>110 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>56</ID>
<type>DE_TO</type>
<position>31,-53.5</position>
<input>
<ID>IN_0</ID>111 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>57</ID>
<type>DE_TO</type>
<position>31,-51.5</position>
<input>
<ID>IN_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>58</ID>
<type>DE_TO</type>
<position>31,-49.5</position>
<input>
<ID>IN_0</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>59</ID>
<type>DE_TO</type>
<position>31,-47.5</position>
<input>
<ID>IN_0</ID>114 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C4</lparam></gate>
<gate>
<ID>60</ID>
<type>DE_TO</type>
<position>31,-45.5</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C5</lparam></gate>
<gate>
<ID>61</ID>
<type>AE_REGISTER8</type>
<position>-7,-19.5</position>
<input>
<ID>IN_0</ID>141 </input>
<input>
<ID>IN_1</ID>146 </input>
<input>
<ID>IN_2</ID>144 </input>
<input>
<ID>IN_3</ID>147 </input>
<input>
<ID>IN_4</ID>140 </input>
<input>
<ID>IN_5</ID>143 </input>
<input>
<ID>IN_6</ID>142 </input>
<input>
<ID>IN_7</ID>145 </input>
<output>
<ID>OUT_0</ID>123 </output>
<output>
<ID>OUT_1</ID>121 </output>
<output>
<ID>OUT_2</ID>116 </output>
<output>
<ID>OUT_3</ID>119 </output>
<output>
<ID>OUT_4</ID>122 </output>
<output>
<ID>OUT_5</ID>120 </output>
<output>
<ID>OUT_6</ID>118 </output>
<output>
<ID>OUT_7</ID>117 </output>
<input>
<ID>clear</ID>174 </input>
<input>
<ID>clock</ID>175 </input>
<input>
<ID>count_enable</ID>173 </input>
<input>
<ID>count_up</ID>173 </input>
<input>
<ID>load</ID>172 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>62</ID>
<type>BW_8X1_BUS_END</type>
<position>-1,-19</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>121 </input>
<input>
<ID>IN_2</ID>116 </input>
<input>
<ID>IN_3</ID>119 </input>
<input>
<ID>IN_4</ID>122 </input>
<input>
<ID>IN_5</ID>120 </input>
<input>
<ID>IN_6</ID>118 </input>
<input>
<ID>IN_7</ID>117 </input>
<input>
<ID>OUT</ID>132 133 134 135 136 137 138 139 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>63</ID>
<type>BW_8X1_BUS_END</type>
<position>14,-19</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>125 </input>
<input>
<ID>IN_2</ID>131 </input>
<input>
<ID>IN_3</ID>124 </input>
<input>
<ID>IN_4</ID>127 </input>
<input>
<ID>IN_5</ID>126 </input>
<input>
<ID>IN_6</ID>129 </input>
<input>
<ID>IN_7</ID>128 </input>
<input>
<ID>OUT</ID>132 133 134 135 136 137 138 139 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>64</ID>
<type>BW_8X1_BUS_END</type>
<position>-13,-19</position>
<input>
<ID>IN_0</ID>141 </input>
<input>
<ID>IN_1</ID>146 </input>
<input>
<ID>IN_2</ID>144 </input>
<input>
<ID>IN_3</ID>147 </input>
<input>
<ID>IN_4</ID>140 </input>
<input>
<ID>IN_5</ID>143 </input>
<input>
<ID>IN_6</ID>142 </input>
<input>
<ID>IN_7</ID>145 </input>
<input>
<ID>OUT</ID>81 82 83 84 85 86 87 88 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>66</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>7,-26</position>
<input>
<ID>ENABLE_0</ID>177 </input>
<input>
<ID>IN_0</ID>148 </input>
<input>
<ID>IN_1</ID>153 </input>
<input>
<ID>IN_2</ID>149 </input>
<input>
<ID>IN_3</ID>151 </input>
<input>
<ID>IN_4</ID>150 </input>
<input>
<ID>IN_5</ID>154 </input>
<input>
<ID>IN_6</ID>152 </input>
<input>
<ID>IN_7</ID>155 </input>
<output>
<ID>OUT_0</ID>156 </output>
<output>
<ID>OUT_1</ID>160 </output>
<output>
<ID>OUT_2</ID>162 </output>
<output>
<ID>OUT_3</ID>158 </output>
<output>
<ID>OUT_4</ID>161 </output>
<output>
<ID>OUT_5</ID>163 </output>
<output>
<ID>OUT_6</ID>159 </output>
<output>
<ID>OUT_7</ID>157 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>67</ID>
<type>BW_8X1_BUS_END</type>
<position>7,-22</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>152 </input>
<input>
<ID>IN_2</ID>154 </input>
<input>
<ID>IN_3</ID>150 </input>
<input>
<ID>IN_4</ID>151 </input>
<input>
<ID>IN_5</ID>149 </input>
<input>
<ID>IN_6</ID>153 </input>
<input>
<ID>IN_7</ID>148 </input>
<input>
<ID>OUT</ID>132 133 134 135 136 137 138 139 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>68</ID>
<type>BW_8X1_BUS_END</type>
<position>7,-30</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>159 </input>
<input>
<ID>IN_2</ID>163 </input>
<input>
<ID>IN_3</ID>161 </input>
<input>
<ID>IN_4</ID>158 </input>
<input>
<ID>IN_5</ID>162 </input>
<input>
<ID>IN_6</ID>160 </input>
<input>
<ID>IN_7</ID>156 </input>
<input>
<ID>OUT</ID>81 82 83 84 85 86 87 88 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>72</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>92,-30</position>
<input>
<ID>ENABLE_0</ID>188 </input>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>109 </input>
<input>
<ID>IN_3</ID>108 </input>
<input>
<ID>IN_4</ID>107 </input>
<input>
<ID>IN_5</ID>106 </input>
<input>
<ID>IN_6</ID>105 </input>
<input>
<ID>IN_7</ID>104 </input>
<output>
<ID>OUT_0</ID>171 </output>
<output>
<ID>OUT_1</ID>170 </output>
<output>
<ID>OUT_2</ID>168 </output>
<output>
<ID>OUT_3</ID>169 </output>
<output>
<ID>OUT_4</ID>164 </output>
<output>
<ID>OUT_5</ID>167 </output>
<output>
<ID>OUT_6</ID>166 </output>
<output>
<ID>OUT_7</ID>165 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>74</ID>
<type>DA_FROM</type>
<position>-14,-11.5</position>
<input>
<ID>IN_0</ID>172 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Counter_load</lparam></gate>
<gate>
<ID>76</ID>
<type>EE_VDD</type>
<position>-7,-9.5</position>
<output>
<ID>OUT_0</ID>173 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>-8,-29.5</position>
<input>
<ID>IN_0</ID>174 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>79</ID>
<type>DA_FROM</type>
<position>-10,-26.5</position>
<input>
<ID>IN_0</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>0.5,-33</position>
<input>
<ID>IN_0</ID>177 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Pass_pointer</lparam></gate>
<gate>
<ID>81</ID>
<type>DA_FROM</type>
<position>59,-4.5</position>
<input>
<ID>IN_0</ID>179 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Pass_addr</lparam></gate>
<gate>
<ID>90</ID>
<type>DE_TO</type>
<position>31,-41.5</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C7</lparam></gate>
<gate>
<ID>92</ID>
<type>DA_FROM</type>
<position>84.5,-30</position>
<input>
<ID>IN_0</ID>188 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Register_store</lparam></gate>
<gate>
<ID>39</ID>
<type>DA_FROM</type>
<position>71.5,-16</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R6</lparam></gate>
<gate>
<ID>103</ID>
<type>DE_TO</type>
<position>-12,-1</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>32</ID>
<type>BB_CLOCK</type>
<position>-20,4.5</position>
<output>
<ID>CLK</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>41</ID>
<type>DA_FROM</type>
<position>76.5,-15</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R7</lparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>100.5,-16</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>54</ID>
<type>DE_TO</type>
<position>105.5,-15</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>65</ID>
<type>DE_TO</type>
<position>106,-32</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>69</ID>
<type>DE_TO</type>
<position>111,-31</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<wire>
<ID>127 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-18.5,16,-18.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_4</name></connection>
<connection>
<GID>63</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>63 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-36,43.5,-36</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<connection>
<GID>20</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>183 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-17.5,35,-14.5</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-17.5,35,-17.5</points>
<connection>
<GID>6</GID>
<name>ENABLE_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>124 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-19.5,16,-19.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_3</name></connection>
<connection>
<GID>63</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>60 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-34,43.5,-34</points>
<connection>
<GID>22</GID>
<name>IN_4</name></connection>
<connection>
<GID>20</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>180 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-29.5,45.5,-27</points>
<connection>
<GID>22</GID>
<name>ENABLE_0</name></connection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-27,49,-27</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>185 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-43.5,18.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_14</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-43.5,29,-43.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-38,43.5,-38</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>186 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-41.5,17.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_15</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-41.5,29,-41.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-37,43.5,-37</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<connection>
<GID>20</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>126 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-17.5,16,-17.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_5</name></connection>
<connection>
<GID>63</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>62 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-35,43.5,-35</points>
<connection>
<GID>22</GID>
<name>IN_3</name></connection>
<connection>
<GID>20</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>128 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-15.5,16,-15.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_7</name></connection>
<connection>
<GID>63</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>64 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-33,43.5,-33</points>
<connection>
<GID>22</GID>
<name>IN_5</name></connection>
<connection>
<GID>20</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>59 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-32,43.5,-32</points>
<connection>
<GID>22</GID>
<name>IN_6</name></connection>
<connection>
<GID>20</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>125 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-21.5,16,-21.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>63</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>61 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-31,43.5,-31</points>
<connection>
<GID>22</GID>
<name>IN_7</name></connection>
<connection>
<GID>20</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>131 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-20.5,16,-20.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_2</name></connection>
<connection>
<GID>63</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>67 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-38,47.5,-38</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>130 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-22.5,16,-22.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>63</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>66 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-37,47.5,-37</points>
<connection>
<GID>22</GID>
<name>OUT_1</name></connection>
<connection>
<GID>24</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>72 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-36,47.5,-36</points>
<connection>
<GID>22</GID>
<name>OUT_2</name></connection>
<connection>
<GID>24</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>129 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-16.5,16,-16.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_6</name></connection>
<connection>
<GID>63</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>65 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-35,47.5,-35</points>
<connection>
<GID>22</GID>
<name>OUT_3</name></connection>
<connection>
<GID>24</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>68 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-34,47.5,-34</points>
<connection>
<GID>22</GID>
<name>OUT_4</name></connection>
<connection>
<GID>24</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>69 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-33,47.5,-33</points>
<connection>
<GID>22</GID>
<name>OUT_5</name></connection>
<connection>
<GID>24</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>71 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-32,47.5,-32</points>
<connection>
<GID>22</GID>
<name>OUT_6</name></connection>
<connection>
<GID>24</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>70 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-31,47.5,-31</points>
<connection>
<GID>22</GID>
<name>OUT_7</name></connection>
<connection>
<GID>24</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>165 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>95.5,-32,95.5,-32</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<connection>
<GID>72</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>166 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>94.5,-32,94.5,-32</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<connection>
<GID>72</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>167 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>93.5,-32,93.5,-32</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<connection>
<GID>72</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>164 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>92.5,-32,92.5,-32</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<connection>
<GID>72</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>169 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>91.5,-32,91.5,-32</points>
<connection>
<GID>70</GID>
<name>IN_4</name></connection>
<connection>
<GID>72</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>168 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>90.5,-32,90.5,-32</points>
<connection>
<GID>70</GID>
<name>IN_5</name></connection>
<connection>
<GID>72</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>170 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>89.5,-32,89.5,-32</points>
<connection>
<GID>70</GID>
<name>IN_6</name></connection>
<connection>
<GID>72</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>171 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>88.5,-32,88.5,-32</points>
<connection>
<GID>70</GID>
<name>IN_7</name></connection>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>81 82 83 84 85 86 87 88 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-39.5,56.5,-27.5</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<intersection>-39.5 1</intersection>
<intersection>-34.5 18</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15,-39.5,98.5,-39.5</points>
<intersection>-15 15</intersection>
<intersection>7 21</intersection>
<intersection>56.5 0</intersection>
<intersection>92 19</intersection>
<intersection>98.5 17</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-15,-39.5,-15,-19</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<intersection>-39.5 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>98.5,-39.5,98.5,-34.5</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>51.5,-34.5,56.5,-34.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>92,-39.5,92,-36</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>-39.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>7,-39.5,7,-32</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>-39.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>28 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-29,32.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>9</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>27 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-29,31.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>9</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>112 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-51.5,22.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_10</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-51.5,29,-51.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49 50 51 52 53 54 55 56 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-34.5,38.5,-16.5</points>
<intersection>-34.5 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-16.5,46.5,-16.5</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-34.5,39.5,-34.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>29 3</intersection>
<intersection>38.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>29,-34.5,29,-33</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>-34.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>113 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-49.5,21.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_11</name></connection>
<intersection>-49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-49.5,29,-49.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-47.5,20.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_12</name></connection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-47.5,29,-47.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-45.5,19.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_13</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-45.5,29,-45.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-29,30.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>9</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>31 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-29,29.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>9</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>29 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-29,28.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>9</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>30 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-29,27.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>9</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>32 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-29,26.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>9</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>25 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-29,25.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>9</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>110 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-55.5,24.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_8</name></connection>
<intersection>-55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-55.5,29,-55.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>111 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-53.5,23.5,-28</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_9</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-53.5,29,-53.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>182 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-15,61.5,-9.5</points>
<connection>
<GID>18</GID>
<name>write_clock</name></connection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>61,-9.5,61.5,-9.5</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-20,51.5,-20</points>
<connection>
<GID>18</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>46 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-19,51.5,-19</points>
<connection>
<GID>18</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>19</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>47 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-18,51.5,-18</points>
<connection>
<GID>18</GID>
<name>ADDRESS_2</name></connection>
<connection>
<GID>19</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>45 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-17,51.5,-17</points>
<connection>
<GID>18</GID>
<name>ADDRESS_3</name></connection>
<connection>
<GID>19</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>48 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-16,51.5,-16</points>
<connection>
<GID>18</GID>
<name>ADDRESS_4</name></connection>
<connection>
<GID>19</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>42 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-15,51.5,-15</points>
<connection>
<GID>18</GID>
<name>ADDRESS_5</name></connection>
<connection>
<GID>19</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>43 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-14,51.5,-14</points>
<connection>
<GID>18</GID>
<name>ADDRESS_6</name></connection>
<connection>
<GID>19</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>44 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-13,51.5,-13</points>
<connection>
<GID>18</GID>
<name>ADDRESS_7</name></connection>
<connection>
<GID>19</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>73 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-23.5,60,-23.5</points>
<connection>
<GID>18</GID>
<name>DATA_IN_0</name></connection>
<connection>
<GID>18</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>77 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-23.5,59,-23.5</points>
<connection>
<GID>18</GID>
<name>DATA_IN_1</name></connection>
<connection>
<GID>18</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>25</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>78 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-23.5,58,-23.5</points>
<connection>
<GID>18</GID>
<name>DATA_IN_2</name></connection>
<connection>
<GID>18</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>25</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>74 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-23.5,57,-23.5</points>
<connection>
<GID>18</GID>
<name>DATA_IN_3</name></connection>
<connection>
<GID>18</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>25</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>79 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-23.5,56,-23.5</points>
<connection>
<GID>18</GID>
<name>DATA_IN_4</name></connection>
<connection>
<GID>18</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>25</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>80 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-23.5,55,-23.5</points>
<connection>
<GID>18</GID>
<name>DATA_IN_5</name></connection>
<connection>
<GID>18</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>25</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>75 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-23.5,54,-23.5</points>
<connection>
<GID>18</GID>
<name>DATA_IN_6</name></connection>
<connection>
<GID>18</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>25</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>76 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-23.5,53,-23.5</points>
<connection>
<GID>18</GID>
<name>DATA_IN_7</name></connection>
<connection>
<GID>18</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>25</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>179 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-17,63,-4.5</points>
<intersection>-17 1</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-17,63,-17</points>
<connection>
<GID>18</GID>
<name>ENABLE_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61,-4.5,63,-4.5</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>181 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-16,62.5,-7</points>
<intersection>-16 1</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-16,62.5,-16</points>
<connection>
<GID>18</GID>
<name>write_enable</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61,-7,62.5,-7</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>184 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-13,82,-12</points>
<connection>
<GID>31</GID>
<name>load</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-12,82,-12</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>187 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-25,82,-24</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<connection>
<GID>31</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>98 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-38,104,-38</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>99 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-37,109,-37</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<connection>
<GID>43</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>100 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-36,104,-36</points>
<connection>
<GID>27</GID>
<name>IN_2</name></connection>
<connection>
<GID>44</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>101 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-35,109,-35</points>
<connection>
<GID>27</GID>
<name>IN_3</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>102 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-34,104,-34</points>
<connection>
<GID>27</GID>
<name>IN_4</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>103 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-33,109,-33</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>102.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>102.5,-33,102.5,-33</points>
<connection>
<GID>27</GID>
<name>IN_5</name></connection>
<intersection>-33 1</intersection></vsegment></shape></wire>
<wire>
<ID>89 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-22,79,-22</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<connection>
<GID>33</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>91 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78.5,-21,79,-21</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<connection>
<GID>34</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>94 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-20,79,-20</points>
<connection>
<GID>31</GID>
<name>IN_2</name></connection>
<connection>
<GID>35</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>92 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78.5,-19,79,-19</points>
<connection>
<GID>31</GID>
<name>IN_3</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>97 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-18,79,-18</points>
<connection>
<GID>31</GID>
<name>IN_4</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>96 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>78.5,-17,79,-17</points>
<connection>
<GID>31</GID>
<name>IN_5</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>104 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87,-22,98.5,-22</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>95.5 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>95.5,-28,95.5,-22</points>
<connection>
<GID>72</GID>
<name>IN_7</name></connection>
<intersection>-22 1</intersection></vsegment></shape></wire>
<wire>
<ID>105 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87,-21,103.5,-21</points>
<connection>
<GID>31</GID>
<name>OUT_1</name></connection>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>94.5 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>94.5,-28,94.5,-21</points>
<connection>
<GID>72</GID>
<name>IN_6</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>106 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87,-20,98.5,-20</points>
<connection>
<GID>31</GID>
<name>OUT_2</name></connection>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>93.5 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>93.5,-28,93.5,-20</points>
<connection>
<GID>72</GID>
<name>IN_5</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>107 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87,-19,103.5,-19</points>
<connection>
<GID>31</GID>
<name>OUT_3</name></connection>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>92.5 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>92.5,-28,92.5,-19</points>
<connection>
<GID>72</GID>
<name>IN_4</name></connection>
<intersection>-19 1</intersection></vsegment></shape></wire>
<wire>
<ID>108 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>87,-18,98.5,-18</points>
<connection>
<GID>31</GID>
<name>OUT_4</name></connection>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>91.5 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>91.5,-28,91.5,-18</points>
<connection>
<GID>72</GID>
<name>IN_3</name></connection>
<intersection>-18 0</intersection></vsegment></shape></wire>
<wire>
<ID>109 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87,-17,103.5,-17</points>
<connection>
<GID>31</GID>
<name>OUT_5</name></connection>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>90.5 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>90.5,-28,90.5,-17</points>
<connection>
<GID>72</GID>
<name>IN_2</name></connection>
<intersection>-17 1</intersection></vsegment></shape></wire>
<wire>
<ID>195 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-15.5,-3.5,-14,-3.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<connection>
<GID>112</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>141 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-11,-22.5,-11,-22.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<connection>
<GID>64</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>146 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-11,-21.5,-11,-21.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<connection>
<GID>64</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>144 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-20.5,-11,-20.5</points>
<connection>
<GID>61</GID>
<name>IN_2</name></connection>
<connection>
<GID>64</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>147 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-19.5,-11,-19.5</points>
<connection>
<GID>61</GID>
<name>IN_3</name></connection>
<connection>
<GID>64</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>140 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-18.5,-11,-18.5</points>
<connection>
<GID>61</GID>
<name>IN_4</name></connection>
<connection>
<GID>64</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>143 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-17.5,-11,-17.5</points>
<connection>
<GID>61</GID>
<name>IN_5</name></connection>
<connection>
<GID>64</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>142 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-16.5,-11,-16.5</points>
<connection>
<GID>61</GID>
<name>IN_6</name></connection>
<connection>
<GID>64</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>145 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-15.5,-11,-15.5</points>
<connection>
<GID>61</GID>
<name>IN_7</name></connection>
<connection>
<GID>64</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>174 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-29.5,-6,-24.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<connection>
<GID>61</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>175 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,-26.5,-8,-24.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<connection>
<GID>61</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>173 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-13.5,-7,-10.5</points>
<connection>
<GID>61</GID>
<name>count_enable</name></connection>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>-13.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-7,-13.5,-6,-13.5</points>
<connection>
<GID>61</GID>
<name>count_up</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>172 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,-13.5,-8,-11.5</points>
<connection>
<GID>61</GID>
<name>load</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,-11.5,-8,-11.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-8 0</intersection></hsegment></shape></wire>
<wire>
<ID>123 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-22.5,-3,-22.5</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<connection>
<GID>62</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>121 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-21.5,-3,-21.5</points>
<connection>
<GID>61</GID>
<name>OUT_1</name></connection>
<connection>
<GID>62</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>116 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-20.5,-3,-20.5</points>
<connection>
<GID>61</GID>
<name>OUT_2</name></connection>
<connection>
<GID>62</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>119 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-19.5,-3,-19.5</points>
<connection>
<GID>61</GID>
<name>OUT_3</name></connection>
<connection>
<GID>62</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>122 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-18.5,-3,-18.5</points>
<connection>
<GID>61</GID>
<name>OUT_4</name></connection>
<connection>
<GID>62</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>120 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-17.5,-3,-17.5</points>
<connection>
<GID>61</GID>
<name>OUT_5</name></connection>
<connection>
<GID>62</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>118 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-16.5,-3,-16.5</points>
<connection>
<GID>61</GID>
<name>OUT_6</name></connection>
<connection>
<GID>62</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>117 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-15.5,-3,-15.5</points>
<connection>
<GID>61</GID>
<name>OUT_7</name></connection>
<connection>
<GID>62</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>132 133 134 135 136 137 138 139 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1,-19,12,-19</points>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>7 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>7,-20,7,-19</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>-19 1</intersection></vsegment></shape></wire>
<wire>
<ID>177 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-33,2.5,-26</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,-26,12,-26</points>
<connection>
<GID>66</GID>
<name>ENABLE_0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>148 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-24,3.5,-24</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<connection>
<GID>67</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>153 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-24,4.5,-24</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<connection>
<GID>67</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>149 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-24,5.5,-24</points>
<connection>
<GID>66</GID>
<name>IN_2</name></connection>
<connection>
<GID>67</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>151 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-24,6.5,-24</points>
<connection>
<GID>66</GID>
<name>IN_3</name></connection>
<connection>
<GID>67</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>150 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-24,7.5,-24</points>
<connection>
<GID>66</GID>
<name>IN_4</name></connection>
<connection>
<GID>67</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>154 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-24,8.5,-24</points>
<connection>
<GID>66</GID>
<name>IN_5</name></connection>
<connection>
<GID>67</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>152 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-24,9.5,-24</points>
<connection>
<GID>66</GID>
<name>IN_6</name></connection>
<connection>
<GID>67</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>155 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-24,10.5,-24</points>
<connection>
<GID>66</GID>
<name>IN_7</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>156 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-28,3.5,-28</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<connection>
<GID>68</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>160 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-28,4.5,-28</points>
<connection>
<GID>66</GID>
<name>OUT_1</name></connection>
<connection>
<GID>68</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>162 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-28,5.5,-28</points>
<connection>
<GID>66</GID>
<name>OUT_2</name></connection>
<connection>
<GID>68</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>158 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-28,6.5,-28</points>
<connection>
<GID>66</GID>
<name>OUT_3</name></connection>
<connection>
<GID>68</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>161 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-28,7.5,-28</points>
<connection>
<GID>66</GID>
<name>OUT_4</name></connection>
<connection>
<GID>68</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>163 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-28,8.5,-28</points>
<connection>
<GID>66</GID>
<name>OUT_5</name></connection>
<connection>
<GID>68</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>159 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-28,9.5,-28</points>
<connection>
<GID>66</GID>
<name>OUT_6</name></connection>
<connection>
<GID>68</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>157 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-28,10.5,-28</points>
<connection>
<GID>66</GID>
<name>OUT_7</name></connection>
<connection>
<GID>68</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>188 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-30,97,-30</points>
<connection>
<GID>72</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>92</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-28,89.5,-16</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>-16 1</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-16,98.5,-16</points>
<connection>
<GID>31</GID>
<name>OUT_6</name></connection>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-28,88.5,-15</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>-15 1</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-15,103.5,-15</points>
<connection>
<GID>31</GID>
<name>OUT_7</name></connection>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,-1,-15,4.5</points>
<intersection>-1 1</intersection>
<intersection>4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15,-1,-14,-1</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>-15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-16,4.5,-15,4.5</points>
<connection>
<GID>32</GID>
<name>CLK</name></connection>
<intersection>-15 0</intersection></hsegment></shape></wire>
<wire>
<ID>11 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-16,79,-16</points>
<connection>
<GID>31</GID>
<name>IN_6</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78.5,-15,79,-15</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<connection>
<GID>31</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>13 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-32,104,-32</points>
<connection>
<GID>27</GID>
<name>IN_6</name></connection>
<connection>
<GID>65</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-31,109,-31</points>
<connection>
<GID>27</GID>
<name>IN_7</name></connection>
<connection>
<GID>69</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-2.07432,5.84775,173.558,-80.0811</PageViewport>
<gate>
<ID>552</ID>
<type>HA_JUNC_2</type>
<position>85.5,-35.5</position>
<input>
<ID>N_in0</ID>592 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>BI_DECODER_4x16</type>
<position>41,-18.5</position>
<input>
<ID>ENABLE</ID>196 </input>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>548 </input>
<input>
<ID>IN_2</ID>547 </input>
<input>
<ID>IN_3</ID>549 </input>
<output>
<ID>OUT_0</ID>565 </output>
<output>
<ID>OUT_1</ID>564 </output>
<output>
<ID>OUT_10</ID>556 </output>
<output>
<ID>OUT_11</ID>555 </output>
<output>
<ID>OUT_12</ID>551 </output>
<output>
<ID>OUT_13</ID>552 </output>
<output>
<ID>OUT_14</ID>550 </output>
<output>
<ID>OUT_15</ID>553 </output>
<output>
<ID>OUT_2</ID>563 </output>
<output>
<ID>OUT_3</ID>562 </output>
<output>
<ID>OUT_4</ID>561 </output>
<output>
<ID>OUT_5</ID>560 </output>
<output>
<ID>OUT_6</ID>558 </output>
<output>
<ID>OUT_7</ID>559 </output>
<output>
<ID>OUT_8</ID>554 </output>
<output>
<ID>OUT_9</ID>557 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>512</ID>
<type>HA_JUNC_2</type>
<position>85.5,-16.5</position>
<input>
<ID>N_in0</ID>557 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>497</ID>
<type>EE_VDD</type>
<position>18,-24</position>
<output>
<ID>OUT_0</ID>541 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>514</ID>
<type>HA_JUNC_2</type>
<position>85.5,-19</position>
<input>
<ID>N_in0</ID>559 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>BA_DECODER_2x4</type>
<position>23,-29.5</position>
<input>
<ID>ENABLE</ID>541 </input>
<input>
<ID>IN_0</ID>540 </input>
<output>
<ID>OUT_0</ID>602 </output>
<output>
<ID>OUT_1</ID>196 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>495</ID>
<type>DA_FROM</type>
<position>17.5,-31</position>
<input>
<ID>IN_0</ID>540 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C4</lparam></gate>
<gate>
<ID>14</ID>
<type>FF_GND</type>
<position>64,-48.5</position>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>516</ID>
<type>HA_JUNC_2</type>
<position>85.5,-21</position>
<input>
<ID>N_in0</ID>560 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AE_OR4</type>
<position>72.5,-54.5</position>
<input>
<ID>IN_0</ID>599 </input>
<input>
<ID>IN_1</ID>597 </input>
<input>
<ID>IN_2</ID>600 </input>
<input>
<ID>IN_3</ID>601 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>502</ID>
<type>DA_FROM</type>
<position>30,-25</position>
<input>
<ID>IN_0</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>503</ID>
<type>DA_FROM</type>
<position>35,-26</position>
<input>
<ID>IN_0</ID>546 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>504</ID>
<type>DA_FROM</type>
<position>30,-23</position>
<input>
<ID>IN_0</ID>549 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>553</ID>
<type>HA_JUNC_2</type>
<position>85.5,-37.5</position>
<input>
<ID>N_in0</ID>590 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>505</ID>
<type>DA_FROM</type>
<position>35,-24</position>
<input>
<ID>IN_0</ID>547 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>520</ID>
<type>HA_JUNC_2</type>
<position>85.5,-25.5</position>
<input>
<ID>N_in0</ID>564 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>506</ID>
<type>HA_JUNC_2</type>
<position>85.5,-10</position>
<input>
<ID>N_in0</ID>553 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>543</ID>
<type>DA_FROM</type>
<position>35,-46</position>
<input>
<ID>IN_0</ID>582 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>507</ID>
<type>HA_JUNC_2</type>
<position>85.5,-11</position>
<input>
<ID>N_in0</ID>550 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>550</ID>
<type>HA_JUNC_2</type>
<position>85.5,-33</position>
<input>
<ID>N_in0</ID>587 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>508</ID>
<type>HA_JUNC_2</type>
<position>85.5,-12</position>
<input>
<ID>N_in0</ID>552 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>557</ID>
<type>HA_JUNC_2</type>
<position>85.5,-44.5</position>
<input>
<ID>N_in0</ID>599 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>509</ID>
<type>HA_JUNC_2</type>
<position>85.5,-13</position>
<input>
<ID>N_in0</ID>551 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>510</ID>
<type>HA_JUNC_2</type>
<position>85.5,-14.5</position>
<input>
<ID>N_in0</ID>555 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>511</ID>
<type>HA_JUNC_2</type>
<position>85.5,-15.5</position>
<input>
<ID>N_in0</ID>556 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>538</ID>
<type>HA_JUNC_2</type>
<position>85.5,-36.5</position>
<input>
<ID>N_in0</ID>593 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>513</ID>
<type>HA_JUNC_2</type>
<position>85.5,-17.5</position>
<input>
<ID>N_in0</ID>554 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>515</ID>
<type>HA_JUNC_2</type>
<position>85.5,-20</position>
<input>
<ID>N_in0</ID>558 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>517</ID>
<type>HA_JUNC_2</type>
<position>85.5,-22</position>
<input>
<ID>N_in0</ID>561 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>518</ID>
<type>HA_JUNC_2</type>
<position>85.5,-23.5</position>
<input>
<ID>N_in0</ID>562 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>519</ID>
<type>HA_JUNC_2</type>
<position>85.5,-24.5</position>
<input>
<ID>N_in0</ID>563 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>DE_TO</type>
<position>59,-58</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Pass_addr</lparam></gate>
<gate>
<ID>521</ID>
<type>HA_JUNC_2</type>
<position>85.5,-26.5</position>
<input>
<ID>N_in0</ID>565 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>539</ID>
<type>BI_DECODER_4x16</type>
<position>41,-38.5</position>
<input>
<ID>ENABLE</ID>602 </input>
<input>
<ID>IN_0</ID>582 </input>
<input>
<ID>IN_1</ID>584 </input>
<input>
<ID>IN_2</ID>583 </input>
<input>
<ID>IN_3</ID>585 </input>
<output>
<ID>OUT_0</ID>601 </output>
<output>
<ID>OUT_1</ID>600 </output>
<output>
<ID>OUT_10</ID>592 </output>
<output>
<ID>OUT_11</ID>591 </output>
<output>
<ID>OUT_12</ID>587 </output>
<output>
<ID>OUT_13</ID>588 </output>
<output>
<ID>OUT_14</ID>586 </output>
<output>
<ID>OUT_15</ID>589 </output>
<output>
<ID>OUT_2</ID>599 </output>
<output>
<ID>OUT_3</ID>598 </output>
<output>
<ID>OUT_4</ID>597 </output>
<output>
<ID>OUT_5</ID>596 </output>
<output>
<ID>OUT_6</ID>594 </output>
<output>
<ID>OUT_7</ID>595 </output>
<output>
<ID>OUT_8</ID>590 </output>
<output>
<ID>OUT_9</ID>593 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>540</ID>
<type>HA_JUNC_2</type>
<position>85.5,-39</position>
<input>
<ID>N_in0</ID>595 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>541</ID>
<type>HA_JUNC_2</type>
<position>85.5,-41</position>
<input>
<ID>N_in0</ID>596 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>542</ID>
<type>DA_FROM</type>
<position>30,-45</position>
<input>
<ID>IN_0</ID>584 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>544</ID>
<type>DA_FROM</type>
<position>30,-43</position>
<input>
<ID>IN_0</ID>585 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>545</ID>
<type>HA_JUNC_2</type>
<position>85.5,-45.5</position>
<input>
<ID>N_in0</ID>600 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>546</ID>
<type>DA_FROM</type>
<position>35,-44</position>
<input>
<ID>IN_0</ID>583 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>547</ID>
<type>HA_JUNC_2</type>
<position>85.5,-30</position>
<input>
<ID>N_in0</ID>589 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>548</ID>
<type>HA_JUNC_2</type>
<position>85.5,-31</position>
<input>
<ID>N_in0</ID>586 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>549</ID>
<type>HA_JUNC_2</type>
<position>85.5,-32</position>
<input>
<ID>N_in0</ID>588 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>551</ID>
<type>HA_JUNC_2</type>
<position>85.5,-34.5</position>
<input>
<ID>N_in0</ID>591 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>554</ID>
<type>HA_JUNC_2</type>
<position>85.5,-40</position>
<input>
<ID>N_in0</ID>594 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>555</ID>
<type>HA_JUNC_2</type>
<position>85.5,-42</position>
<input>
<ID>N_in0</ID>597 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>556</ID>
<type>HA_JUNC_2</type>
<position>85.5,-43.5</position>
<input>
<ID>N_in0</ID>598 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>558</ID>
<type>HA_JUNC_2</type>
<position>85.5,-46.5</position>
<input>
<ID>N_in0</ID>601 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>560</ID>
<type>DE_TO</type>
<position>47.5,-49.5</position>
<input>
<ID>IN_0</ID>598 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Counter_load</lparam></gate>
<gate>
<ID>1</ID>
<type>DE_TO</type>
<position>51,-55.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Pass_value</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_OR2</type>
<position>51,-50.5</position>
<input>
<ID>IN_0</ID>564 </input>
<input>
<ID>IN_1</ID>600 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>DM_NOR8</type>
<position>59,-50.5</position>
<input>
<ID>IN_0</ID>599 </input>
<input>
<ID>IN_1</ID>601 </input>
<input>
<ID>IN_2</ID>595 </input>
<input>
<ID>IN_3</ID>594 </input>
<input>
<ID>IN_4</ID>600 </input>
<input>
<ID>IN_5</ID>564 </input>
<input>
<ID>IN_6</ID>597 </input>
<input>
<ID>IN_7</ID>596 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>15</ID>
<type>DE_TO</type>
<position>66.5,-51</position>
<input>
<ID>IN_0</ID>599 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Pass_pointer</lparam></gate>
<gate>
<ID>17</ID>
<type>DE_TO</type>
<position>72.5,-60.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID write</lparam></gate>
<gate>
<ID>26</ID>
<type>DE_TO</type>
<position>79,-51</position>
<input>
<ID>IN_0</ID>601 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Register_store</lparam></gate>
<wire>
<ID>565 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-26.5,84.5,-26.5</points>
<connection>
<GID>521</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-26.5,44,-26</points>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection>
<intersection>-26.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>549 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-23,38,-23</points>
<connection>
<GID>504</GID>
<name>IN_0</name></connection>
<connection>
<GID>114</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>541 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-28,18,-25</points>
<connection>
<GID>497</GID>
<name>OUT_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-28,20,-28</points>
<connection>
<GID>120</GID>
<name>ENABLE</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>557 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-16.5,84.5,-16.5</points>
<connection>
<GID>512</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-17,44,-16.5</points>
<connection>
<GID>114</GID>
<name>OUT_9</name></connection>
<intersection>-16.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>592 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-35.5,84.5,-35.5</points>
<connection>
<GID>552</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-36,44,-35.5</points>
<connection>
<GID>539</GID>
<name>OUT_10</name></connection>
<intersection>-35.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>590 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-37.5,84.5,-37.5</points>
<connection>
<GID>553</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-38,44,-37.5</points>
<connection>
<GID>539</GID>
<name>OUT_8</name></connection>
<intersection>-37.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>196 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-30,33.5,-11</points>
<intersection>-30 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-11,38,-11</points>
<connection>
<GID>114</GID>
<name>ENABLE</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-30,33.5,-30</points>
<connection>
<GID>120</GID>
<name>OUT_1</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>546 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-26,38,-26</points>
<connection>
<GID>503</GID>
<name>IN_0</name></connection>
<connection>
<GID>114</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>548 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-25,38,-25</points>
<connection>
<GID>502</GID>
<name>IN_0</name></connection>
<connection>
<GID>114</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>547 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-24,38,-24</points>
<connection>
<GID>505</GID>
<name>IN_0</name></connection>
<connection>
<GID>114</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>564 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-25.5,84.5,-25.5</points>
<connection>
<GID>520</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection>
<intersection>52 8</intersection>
<intersection>56.5 10</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-25.5,44,-25</points>
<connection>
<GID>114</GID>
<name>OUT_1</name></connection>
<intersection>-25.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>52,-47.5,52,-25.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>-25.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>56.5,-47.5,56.5,-25.5</points>
<connection>
<GID>12</GID>
<name>IN_5</name></connection>
<intersection>-25.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>556 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-15.5,84.5,-15.5</points>
<connection>
<GID>511</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-16,44,-15.5</points>
<connection>
<GID>114</GID>
<name>OUT_10</name></connection>
<intersection>-15.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>555 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-14.5,84.5,-14.5</points>
<connection>
<GID>510</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-15,44,-14.5</points>
<connection>
<GID>114</GID>
<name>OUT_11</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>551 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-13,84.5,-13</points>
<connection>
<GID>509</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-14,44,-13</points>
<connection>
<GID>114</GID>
<name>OUT_12</name></connection>
<intersection>-13 1</intersection></vsegment></shape></wire>
<wire>
<ID>552 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-12,84.5,-12</points>
<connection>
<GID>508</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-13,44,-12</points>
<connection>
<GID>114</GID>
<name>OUT_13</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire>
<wire>
<ID>550 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-11,84.5,-11</points>
<connection>
<GID>507</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-12,44,-11</points>
<connection>
<GID>114</GID>
<name>OUT_14</name></connection>
<intersection>-11 1</intersection></vsegment></shape></wire>
<wire>
<ID>553 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-10,84.5,-10</points>
<connection>
<GID>506</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-11,44,-10</points>
<connection>
<GID>114</GID>
<name>OUT_15</name></connection>
<intersection>-10 1</intersection></vsegment></shape></wire>
<wire>
<ID>563 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-24.5,84.5,-24.5</points>
<connection>
<GID>519</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-24.5,44,-24</points>
<connection>
<GID>114</GID>
<name>OUT_2</name></connection>
<intersection>-24.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>562 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-23.5,84.5,-23.5</points>
<connection>
<GID>518</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-23.5,44,-23</points>
<connection>
<GID>114</GID>
<name>OUT_3</name></connection>
<intersection>-23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>561 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-22,84.5,-22</points>
<connection>
<GID>517</GID>
<name>N_in0</name></connection>
<connection>
<GID>114</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>560 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-21,84.5,-21</points>
<connection>
<GID>516</GID>
<name>N_in0</name></connection>
<connection>
<GID>114</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>558 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-20,84.5,-20</points>
<connection>
<GID>515</GID>
<name>N_in0</name></connection>
<connection>
<GID>114</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>559 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-19,84.5,-19</points>
<connection>
<GID>514</GID>
<name>N_in0</name></connection>
<connection>
<GID>114</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>554 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-17.5,84.5,-17.5</points>
<connection>
<GID>513</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-18,44,-17.5</points>
<connection>
<GID>114</GID>
<name>OUT_8</name></connection>
<intersection>-17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>540 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-31,20,-31</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<connection>
<GID>120</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>602 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-31,38,-31</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<connection>
<GID>539</GID>
<name>ENABLE</name></connection></hsegment></shape></wire>
<wire>
<ID>582 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-46,38,-46</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<connection>
<GID>543</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>587 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-33,84.5,-33</points>
<connection>
<GID>550</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-34,44,-33</points>
<connection>
<GID>539</GID>
<name>OUT_12</name></connection>
<intersection>-33 1</intersection></vsegment></shape></wire>
<wire>
<ID>599 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-44.5,84.5,-44.5</points>
<connection>
<GID>557</GID>
<name>N_in0</name></connection>
<intersection>44 11</intersection>
<intersection>62.5 14</intersection>
<intersection>66.5 12</intersection>
<intersection>75.5 16</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>44,-44.5,44,-44</points>
<connection>
<GID>539</GID>
<name>OUT_2</name></connection>
<intersection>-44.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>66.5,-49,66.5,-44.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-44.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>62.5,-47.5,62.5,-44.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-44.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>75.5,-51.5,75.5,-44.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>-44.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>593 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-36.5,84.5,-36.5</points>
<connection>
<GID>538</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-37,44,-36.5</points>
<connection>
<GID>539</GID>
<name>OUT_9</name></connection>
<intersection>-36.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>584 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-45,38,-45</points>
<connection>
<GID>542</GID>
<name>IN_0</name></connection>
<connection>
<GID>539</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>9 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-58.5,72.5,-58.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<connection>
<GID>17</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>583 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-44,38,-44</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<connection>
<GID>539</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>585 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-43,38,-43</points>
<connection>
<GID>544</GID>
<name>IN_0</name></connection>
<connection>
<GID>539</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>601 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-46.5,84.5,-46.5</points>
<connection>
<GID>558</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection>
<intersection>61.5 10</intersection>
<intersection>69.5 8</intersection>
<intersection>79 9</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-46.5,44,-46</points>
<connection>
<GID>539</GID>
<name>OUT_0</name></connection>
<intersection>-46.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>69.5,-51.5,69.5,-46.5</points>
<connection>
<GID>29</GID>
<name>IN_3</name></connection>
<intersection>-46.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>79,-49,79,-46.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-46.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>61.5,-47.5,61.5,-46.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>-46.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>600 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-45.5,84.5,-45.5</points>
<connection>
<GID>545</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection>
<intersection>50 8</intersection>
<intersection>55.5 9</intersection>
<intersection>71.5 13</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-45.5,44,-45</points>
<connection>
<GID>539</GID>
<name>OUT_1</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>50,-47.5,50,-45.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>55.5,-47.5,55.5,-45.5</points>
<connection>
<GID>12</GID>
<name>IN_4</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>71.5,-51.5,71.5,-45.5</points>
<connection>
<GID>29</GID>
<name>IN_2</name></connection>
<intersection>-45.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>591 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-34.5,84.5,-34.5</points>
<connection>
<GID>551</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-35,44,-34.5</points>
<connection>
<GID>539</GID>
<name>OUT_11</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>588 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-32,84.5,-32</points>
<connection>
<GID>549</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-33,44,-32</points>
<connection>
<GID>539</GID>
<name>OUT_13</name></connection>
<intersection>-32 1</intersection></vsegment></shape></wire>
<wire>
<ID>586 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-31,84.5,-31</points>
<connection>
<GID>548</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-32,44,-31</points>
<connection>
<GID>539</GID>
<name>OUT_14</name></connection>
<intersection>-31 1</intersection></vsegment></shape></wire>
<wire>
<ID>589 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-30,84.5,-30</points>
<connection>
<GID>547</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-31,44,-30</points>
<connection>
<GID>539</GID>
<name>OUT_15</name></connection>
<intersection>-30 1</intersection></vsegment></shape></wire>
<wire>
<ID>598 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-43.5,84.5,-43.5</points>
<connection>
<GID>556</GID>
<name>N_in0</name></connection>
<intersection>44 7</intersection>
<intersection>47.5 8</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>44,-43.5,44,-43</points>
<connection>
<GID>539</GID>
<name>OUT_3</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>47.5,-47.5,47.5,-43.5</points>
<connection>
<GID>560</GID>
<name>IN_0</name></connection>
<intersection>-43.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-56,59,-54.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>-54.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>59,-54.5,59,-54.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>597 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-42,84.5,-42</points>
<connection>
<GID>555</GID>
<name>N_in0</name></connection>
<connection>
<GID>539</GID>
<name>OUT_4</name></connection>
<intersection>57.5 2</intersection>
<intersection>73.5 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57.5,-47.5,57.5,-42</points>
<connection>
<GID>12</GID>
<name>IN_6</name></connection>
<intersection>-42 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>73.5,-51.5,73.5,-42</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>-42 1</intersection></vsegment></shape></wire>
<wire>
<ID>596 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-41,84.5,-41</points>
<connection>
<GID>541</GID>
<name>N_in0</name></connection>
<connection>
<GID>539</GID>
<name>OUT_5</name></connection>
<intersection>58.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>58.5,-47.5,58.5,-41</points>
<connection>
<GID>12</GID>
<name>IN_7</name></connection>
<intersection>-41 1</intersection></vsegment></shape></wire>
<wire>
<ID>594 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-40,84.5,-40</points>
<connection>
<GID>554</GID>
<name>N_in0</name></connection>
<connection>
<GID>539</GID>
<name>OUT_6</name></connection>
<intersection>59.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>59.5,-47.5,59.5,-40</points>
<connection>
<GID>12</GID>
<name>IN_3</name></connection>
<intersection>-40 1</intersection></vsegment></shape></wire>
<wire>
<ID>595 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-39,84.5,-39</points>
<connection>
<GID>540</GID>
<name>N_in0</name></connection>
<connection>
<GID>539</GID>
<name>OUT_7</name></connection>
<intersection>60.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>60.5,-47.5,60.5,-39</points>
<connection>
<GID>12</GID>
<name>IN_2</name></connection>
<intersection>-39 1</intersection></vsegment></shape></wire>
<wire>
<ID>1 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-53.5,51,-53.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-53.5,51,-53.5</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-53.3179,-27.1114,162.597,-132.749</PageViewport>
<gate>
<ID>185</ID>
<type>DA_FROM</type>
<position>-2.5,-23.5</position>
<input>
<ID>IN_0</ID>259 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>121</ID>
<type>DA_FROM</type>
<position>28,13.5</position>
<input>
<ID>IN_0</ID>270 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>129</ID>
<type>DA_FROM</type>
<position>37.5,-25</position>
<input>
<ID>IN_0</ID>415 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>282</ID>
<type>DA_FROM</type>
<position>48.5,-26</position>
<input>
<ID>IN_0</ID>416 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>122</ID>
<type>DA_FROM</type>
<position>-4.5,-23.5</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>481</ID>
<type>DA_FROM</type>
<position>81,-31</position>
<input>
<ID>IN_0</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR5</lparam></gate>
<gate>
<ID>123</ID>
<type>DA_FROM</type>
<position>47.5,-69</position>
<input>
<ID>IN_0</ID>432 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND2</lparam></gate>
<gate>
<ID>124</ID>
<type>DA_FROM</type>
<position>28,15.5</position>
<input>
<ID>IN_0</ID>267 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>475</ID>
<type>DE_TO</type>
<position>103,-32.5</position>
<input>
<ID>IN_0</ID>480 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R5</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>19.5,4</position>
<input>
<ID>IN_0</ID>204 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>485</ID>
<type>DA_FROM</type>
<position>70.5,-58</position>
<input>
<ID>IN_0</ID>508 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>52.5,-57</position>
<input>
<ID>IN_0</ID>421 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>127</ID>
<type>DE_TO</type>
<position>59.5,2</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0</lparam></gate>
<gate>
<ID>128</ID>
<type>DA_FROM</type>
<position>-0.5,-23.5</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>130</ID>
<type>AM_MUX_16x1</type>
<position>54,2</position>
<input>
<ID>IN_0</ID>267 </input>
<input>
<ID>IN_1</ID>267 </input>
<input>
<ID>IN_10</ID>370 </input>
<input>
<ID>IN_11</ID>399 </input>
<input>
<ID>IN_12</ID>397 </input>
<input>
<ID>IN_13</ID>398 </input>
<input>
<ID>IN_14</ID>396 </input>
<input>
<ID>IN_15</ID>395 </input>
<input>
<ID>IN_2</ID>268 </input>
<input>
<ID>IN_3</ID>269 </input>
<input>
<ID>IN_4</ID>271 </input>
<input>
<ID>IN_5</ID>272 </input>
<input>
<ID>IN_6</ID>295 </input>
<input>
<ID>IN_7</ID>295 </input>
<input>
<ID>IN_8</ID>368 </input>
<input>
<ID>IN_9</ID>369 </input>
<output>
<ID>OUT</ID>198 </output>
<input>
<ID>SEL_0</ID>202 </input>
<input>
<ID>SEL_1</ID>201 </input>
<input>
<ID>SEL_2</ID>199 </input>
<input>
<ID>SEL_3</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>292</ID>
<type>AA_AND2</type>
<position>-40,-21</position>
<input>
<ID>IN_0</ID>315 </input>
<input>
<ID>IN_1</ID>314 </input>
<output>
<ID>OUT</ID>316 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>15.5,4</position>
<input>
<ID>IN_0</ID>206 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>47.5,-65</position>
<input>
<ID>IN_0</ID>437 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>286</ID>
<type>DA_FROM</type>
<position>-45,-18</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>133</ID>
<type>DA_FROM</type>
<position>55.5,14.5</position>
<input>
<ID>IN_0</ID>202 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>134</ID>
<type>DA_FROM</type>
<position>10.5,4</position>
<input>
<ID>IN_0</ID>208 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>280</ID>
<type>AA_AND2</type>
<position>-40,-17</position>
<input>
<ID>IN_0</ID>312 </input>
<input>
<ID>IN_1</ID>311 </input>
<output>
<ID>OUT</ID>313 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>38,-73</position>
<input>
<ID>IN_0</ID>429 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum2</lparam></gate>
<gate>
<ID>136</ID>
<type>DA_FROM</type>
<position>54.5,19.5</position>
<input>
<ID>IN_0</ID>201 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>290</ID>
<type>DA_FROM</type>
<position>5,-108</position>
<input>
<ID>IN_0</ID>377 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>137</ID>
<type>DA_FROM</type>
<position>53.5,14.5</position>
<input>
<ID>IN_0</ID>199 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>138</ID>
<type>DA_FROM</type>
<position>54.5,-57</position>
<input>
<ID>IN_0</ID>424 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>300</ID>
<type>DA_FROM</type>
<position>-45,-60</position>
<input>
<ID>IN_0</ID>334 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>139</ID>
<type>DA_FROM</type>
<position>52.5,19.5</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>140</ID>
<type>DA_FROM</type>
<position>-13.5,-28.5</position>
<input>
<ID>IN_0</ID>239 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>294</ID>
<type>DA_FROM</type>
<position>27,-58</position>
<input>
<ID>IN_0</ID>428 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>141</ID>
<type>DA_FROM</type>
<position>-2.5,4</position>
<input>
<ID>IN_0</ID>214 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>142</ID>
<type>DA_FROM</type>
<position>38,-70.5</position>
<input>
<ID>IN_0</ID>431 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec2</lparam></gate>
<gate>
<ID>288</ID>
<type>DA_FROM</type>
<position>36.5,-62</position>
<input>
<ID>IN_0</ID>435 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>143</ID>
<type>DA_FROM</type>
<position>-4.5,4</position>
<input>
<ID>IN_0</ID>215 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>144</ID>
<type>DE_TO</type>
<position>-13,-43</position>
<input>
<ID>IN_0</ID>248 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID UF</lparam></gate>
<gate>
<ID>298</ID>
<type>DE_TO</type>
<position>-35,-21</position>
<input>
<ID>IN_0</ID>316 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND6</lparam></gate>
<gate>
<ID>145</ID>
<type>DA_FROM</type>
<position>-7.5,4</position>
<input>
<ID>IN_0</ID>216 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>146</ID>
<type>DA_FROM</type>
<position>-9.5,4</position>
<input>
<ID>IN_0</ID>217 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>308</ID>
<type>DA_FROM</type>
<position>80,-64</position>
<input>
<ID>IN_0</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>147</ID>
<type>DA_FROM</type>
<position>-11.5,4</position>
<input>
<ID>IN_0</ID>218 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>148</ID>
<type>DE_TO</type>
<position>8,-42.5</position>
<input>
<ID>IN_0</ID>243 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff3</lparam></gate>
<gate>
<ID>302</ID>
<type>AM_MUX_16x1</type>
<position>53,-105</position>
<input>
<ID>IN_0</ID>445 </input>
<input>
<ID>IN_1</ID>445 </input>
<input>
<ID>IN_10</ID>454 </input>
<input>
<ID>IN_11</ID>459 </input>
<input>
<ID>IN_12</ID>457 </input>
<input>
<ID>IN_13</ID>458 </input>
<input>
<ID>IN_14</ID>456 </input>
<input>
<ID>IN_15</ID>455 </input>
<input>
<ID>IN_2</ID>446 </input>
<input>
<ID>IN_3</ID>447 </input>
<input>
<ID>IN_4</ID>449 </input>
<input>
<ID>IN_5</ID>450 </input>
<input>
<ID>IN_6</ID>451 </input>
<input>
<ID>IN_7</ID>451 </input>
<input>
<ID>IN_8</ID>452 </input>
<input>
<ID>IN_9</ID>453 </input>
<output>
<ID>OUT</ID>440 </output>
<input>
<ID>SEL_0</ID>444 </input>
<input>
<ID>SEL_1</ID>443 </input>
<input>
<ID>SEL_2</ID>441 </input>
<input>
<ID>SEL_3</ID>442 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>149</ID>
<type>DA_FROM</type>
<position>-13.5,4</position>
<input>
<ID>IN_0</ID>219 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>150</ID>
<type>DA_FROM</type>
<position>-9.5,-28.5</position>
<input>
<ID>IN_0</ID>237 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>296</ID>
<type>DA_FROM</type>
<position>-45,-22</position>
<input>
<ID>IN_0</ID>314 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>151</ID>
<type>DE_TO</type>
<position>14,-10</position>
<input>
<ID>IN_0</ID>220 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum0</lparam></gate>
<gate>
<ID>152</ID>
<type>DE_TO</type>
<position>12,-10</position>
<input>
<ID>IN_0</ID>221 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum1</lparam></gate>
<gate>
<ID>306</ID>
<type>DA_FROM</type>
<position>-45,-26</position>
<input>
<ID>IN_0</ID>317 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>153</ID>
<type>DE_TO</type>
<position>-9.5,-42.5</position>
<input>
<ID>IN_0</ID>247 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff7</lparam></gate>
<gate>
<ID>154</ID>
<type>DE_TO</type>
<position>10,-10</position>
<input>
<ID>IN_0</ID>222 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum2</lparam></gate>
<gate>
<ID>316</ID>
<type>DA_FROM</type>
<position>81,9.5</position>
<input>
<ID>IN_0</ID>475 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>155</ID>
<type>DE_TO</type>
<position>8,-10</position>
<input>
<ID>IN_0</ID>223 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum3</lparam></gate>
<gate>
<ID>156</ID>
<type>DE_TO</type>
<position>-3.5,-10</position>
<input>
<ID>IN_0</ID>224 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum4</lparam></gate>
<gate>
<ID>310</ID>
<type>DA_FROM</type>
<position>81,5.5</position>
<input>
<ID>IN_0</ID>479 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>157</ID>
<type>DE_TO</type>
<position>-5.5,-10</position>
<input>
<ID>IN_0</ID>225 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum5</lparam></gate>
<gate>
<ID>158</ID>
<type>DE_TO</type>
<position>-7.5,-10</position>
<input>
<ID>IN_0</ID>226 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum6</lparam></gate>
<gate>
<ID>304</ID>
<type>DA_FROM</type>
<position>-45,-24</position>
<input>
<ID>IN_0</ID>318 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>159</ID>
<type>DE_TO</type>
<position>-9.5,-10</position>
<input>
<ID>IN_0</ID>227 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum7</lparam></gate>
<gate>
<ID>160</ID>
<type>DE_TO</type>
<position>-5.5,-42.5</position>
<input>
<ID>IN_0</ID>245 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff5</lparam></gate>
<gate>
<ID>314</ID>
<type>DA_FROM</type>
<position>-45,-36</position>
<input>
<ID>IN_0</ID>322 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>161</ID>
<type>FF_GND</type>
<position>20,-3.5</position>
<output>
<ID>OUT_0</ID>228 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>162</ID>
<type>DE_TO</type>
<position>-13,-10.5</position>
<input>
<ID>IN_0</ID>229 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID OV</lparam></gate>
<gate>
<ID>163</ID>
<type>DE_TO</type>
<position>-15,-10.5</position>
<input>
<ID>IN_0</ID>230 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Sum8</lparam></gate>
<gate>
<ID>164</ID>
<type>DA_FROM</type>
<position>-7.5,-28.5</position>
<input>
<ID>IN_0</ID>236 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_FROM</type>
<position>-11.5,-28.5</position>
<input>
<ID>IN_0</ID>238 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>318</ID>
<type>DA_FROM</type>
<position>-45,-40</position>
<input>
<ID>IN_0</ID>325 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>166</ID>
<type>DE_TO</type>
<position>14,-42.5</position>
<input>
<ID>IN_0</ID>240 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff0</lparam></gate>
<gate>
<ID>167</ID>
<type>DA_FROM</type>
<position>-0.5,4</position>
<input>
<ID>IN_0</ID>213 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>312</ID>
<type>DA_FROM</type>
<position>-45,-34</position>
<input>
<ID>IN_0</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>168</ID>
<type>DE_TO</type>
<position>12,-42.5</position>
<input>
<ID>IN_0</ID>241 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff1</lparam></gate>
<gate>
<ID>169</ID>
<type>DE_TO</type>
<position>10,-42.5</position>
<input>
<ID>IN_0</ID>242 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff2</lparam></gate>
<gate>
<ID>170</ID>
<type>DE_TO</type>
<position>-3.5,-42.5</position>
<input>
<ID>IN_0</ID>244 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff4</lparam></gate>
<gate>
<ID>171</ID>
<type>DE_TO</type>
<position>-7.5,-42.5</position>
<input>
<ID>IN_0</ID>246 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff6</lparam></gate>
<gate>
<ID>172</ID>
<type>DE_TO</type>
<position>-15,-43</position>
<input>
<ID>IN_0</ID>249 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Diff8</lparam></gate>
<gate>
<ID>173</ID>
<type>AE_FULLADDER_4BIT</type>
<position>11,-35.5</position>
<input>
<ID>IN_0</ID>232 </input>
<input>
<ID>IN_1</ID>233 </input>
<input>
<ID>IN_2</ID>234 </input>
<input>
<ID>IN_3</ID>235 </input>
<input>
<ID>IN_B_0</ID>253 </input>
<input>
<ID>IN_B_1</ID>251 </input>
<input>
<ID>IN_B_2</ID>252 </input>
<input>
<ID>IN_B_3</ID>250 </input>
<output>
<ID>OUT_0</ID>240 </output>
<output>
<ID>OUT_1</ID>241 </output>
<output>
<ID>OUT_2</ID>242 </output>
<output>
<ID>OUT_3</ID>243 </output>
<input>
<ID>carry_in</ID>266 </input>
<output>
<ID>carry_out</ID>231 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>174</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-6.5,-35.5</position>
<input>
<ID>IN_0</ID>236 </input>
<input>
<ID>IN_1</ID>237 </input>
<input>
<ID>IN_2</ID>238 </input>
<input>
<ID>IN_3</ID>239 </input>
<input>
<ID>IN_B_0</ID>262 </input>
<input>
<ID>IN_B_1</ID>263 </input>
<input>
<ID>IN_B_2</ID>264 </input>
<input>
<ID>IN_B_3</ID>265 </input>
<output>
<ID>OUT_0</ID>244 </output>
<output>
<ID>OUT_1</ID>245 </output>
<output>
<ID>OUT_2</ID>246 </output>
<output>
<ID>OUT_3</ID>247 </output>
<input>
<ID>carry_in</ID>231 </input>
<output>
<ID>carry_out</ID>249 </output>
<output>
<ID>overflow</ID>248 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>175</ID>
<type>DA_FROM</type>
<position>19,-23.5</position>
<input>
<ID>IN_0</ID>256 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>176</ID>
<type>DA_FROM</type>
<position>17,-23.5</position>
<input>
<ID>IN_0</ID>257 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>177</ID>
<type>DA_FROM</type>
<position>15,-23.5</position>
<input>
<ID>IN_0</ID>255 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>178</ID>
<type>DA_FROM</type>
<position>13,-23.5</position>
<input>
<ID>IN_0</ID>254 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>179</ID>
<type>DA_FROM</type>
<position>10.5,-28.5</position>
<input>
<ID>IN_0</ID>232 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>180</ID>
<type>DA_FROM</type>
<position>8.5,-28.5</position>
<input>
<ID>IN_0</ID>233 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>181</ID>
<type>DA_FROM</type>
<position>6.5,-28.5</position>
<input>
<ID>IN_0</ID>234 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>182</ID>
<type>DA_FROM</type>
<position>4.5,-28.5</position>
<input>
<ID>IN_0</ID>235 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>183</ID>
<type>AI_INVERTER_4BIT</type>
<position>14.5,-29</position>
<input>
<ID>IN_0</ID>254 </input>
<input>
<ID>IN_1</ID>255 </input>
<input>
<ID>IN_2</ID>257 </input>
<input>
<ID>IN_3</ID>256 </input>
<output>
<ID>OUT_0</ID>250 </output>
<output>
<ID>OUT_1</ID>252 </output>
<output>
<ID>OUT_2</ID>251 </output>
<output>
<ID>OUT_3</ID>253 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>184</ID>
<type>DA_FROM</type>
<position>1.5,-23.5</position>
<input>
<ID>IN_0</ID>260 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>186</ID>
<type>AI_INVERTER_4BIT</type>
<position>-3,-29</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>259 </input>
<input>
<ID>IN_2</ID>261 </input>
<input>
<ID>IN_3</ID>260 </input>
<output>
<ID>OUT_0</ID>265 </output>
<output>
<ID>OUT_1</ID>264 </output>
<output>
<ID>OUT_2</ID>263 </output>
<output>
<ID>OUT_3</ID>262 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>187</ID>
<type>EE_VDD</type>
<position>20,-32.5</position>
<output>
<ID>OUT_0</ID>266 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_LABEL</type>
<position>-6.5,16</position>
<gparam>LABEL_TEXT ALU</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>189</ID>
<type>AE_FULLADDER_4BIT</type>
<position>11,-3</position>
<input>
<ID>IN_0</ID>208 </input>
<input>
<ID>IN_1</ID>209 </input>
<input>
<ID>IN_2</ID>210 </input>
<input>
<ID>IN_3</ID>211 </input>
<input>
<ID>IN_B_0</ID>204 </input>
<input>
<ID>IN_B_1</ID>205 </input>
<input>
<ID>IN_B_2</ID>206 </input>
<input>
<ID>IN_B_3</ID>207 </input>
<output>
<ID>OUT_0</ID>220 </output>
<output>
<ID>OUT_1</ID>221 </output>
<output>
<ID>OUT_2</ID>222 </output>
<output>
<ID>OUT_3</ID>223 </output>
<input>
<ID>carry_in</ID>228 </input>
<output>
<ID>carry_out</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>190</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-6.5,-3</position>
<input>
<ID>IN_0</ID>216 </input>
<input>
<ID>IN_1</ID>217 </input>
<input>
<ID>IN_2</ID>218 </input>
<input>
<ID>IN_3</ID>219 </input>
<input>
<ID>IN_B_0</ID>212 </input>
<input>
<ID>IN_B_1</ID>213 </input>
<input>
<ID>IN_B_2</ID>214 </input>
<input>
<ID>IN_B_3</ID>215 </input>
<output>
<ID>OUT_0</ID>224 </output>
<output>
<ID>OUT_1</ID>225 </output>
<output>
<ID>OUT_2</ID>226 </output>
<output>
<ID>OUT_3</ID>227 </output>
<input>
<ID>carry_in</ID>203 </input>
<output>
<ID>carry_out</ID>230 </output>
<output>
<ID>overflow</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>191</ID>
<type>DA_FROM</type>
<position>17.5,4</position>
<input>
<ID>IN_0</ID>205 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>192</ID>
<type>DA_FROM</type>
<position>13,4</position>
<input>
<ID>IN_0</ID>207 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>193</ID>
<type>DA_FROM</type>
<position>8.5,4</position>
<input>
<ID>IN_0</ID>209 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>346</ID>
<type>DE_TO</type>
<position>-35,-33</position>
<input>
<ID>IN_0</ID>336 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR0</lparam></gate>
<gate>
<ID>194</ID>
<type>DA_FROM</type>
<position>6.5,4</position>
<input>
<ID>IN_0</ID>210 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>195</ID>
<type>DA_FROM</type>
<position>4.5,4</position>
<input>
<ID>IN_0</ID>211 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>356</ID>
<type>DA_FROM</type>
<position>91,-67</position>
<input>
<ID>IN_0</ID>514 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR6</lparam></gate>
<gate>
<ID>196</ID>
<type>DA_FROM</type>
<position>1.5,4</position>
<input>
<ID>IN_0</ID>212 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>197</ID>
<type>DE_TO</type>
<position>-35,-53</position>
<input>
<ID>IN_0</ID>341 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR5</lparam></gate>
<gate>
<ID>350</ID>
<type>DA_FROM</type>
<position>97,-52</position>
<input>
<ID>IN_0</ID>503 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>198</ID>
<type>AE_SMALL_INVERTER</type>
<position>43,-3.5</position>
<input>
<ID>IN_0</ID>267 </input>
<output>
<ID>OUT_0</ID>268 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>199</ID>
<type>AE_SMALL_INVERTER</type>
<position>47.5,-2.5</position>
<input>
<ID>IN_0</ID>270 </input>
<output>
<ID>OUT_0</ID>269 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>344</ID>
<type>DA_FROM</type>
<position>70.5,-56</position>
<input>
<ID>IN_0</ID>505 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>200</ID>
<type>DA_FROM</type>
<position>-45,-80</position>
<input>
<ID>IN_0</ID>349 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>201</ID>
<type>DA_FROM</type>
<position>39,-1.5</position>
<input>
<ID>IN_0</ID>271 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum0</lparam></gate>
<gate>
<ID>354</ID>
<type>DE_TO</type>
<position>-35,-49</position>
<input>
<ID>IN_0</ID>340 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR4</lparam></gate>
<gate>
<ID>202</ID>
<type>DA_FROM</type>
<position>-45,-70</position>
<input>
<ID>IN_0</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>203</ID>
<type>DA_FROM</type>
<position>28.5,-0.5</position>
<input>
<ID>IN_0</ID>272 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff0</lparam></gate>
<gate>
<ID>364</ID>
<type>DA_FROM</type>
<position>-45,-68</position>
<input>
<ID>IN_0</ID>345 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>204</ID>
<type>DA_FROM</type>
<position>-45,-76</position>
<input>
<ID>IN_0</ID>346 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>205</ID>
<type>DA_FROM</type>
<position>10.5,-59.5</position>
<input>
<ID>IN_0</ID>274 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>358</ID>
<type>DA_FROM</type>
<position>-45,-86</position>
<input>
<ID>IN_0</ID>353 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>206</ID>
<type>DA_FROM</type>
<position>-7.5,-59.5</position>
<input>
<ID>IN_0</ID>278 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>207</ID>
<type>DA_FROM</type>
<position>-45,-88</position>
<input>
<ID>IN_0</ID>352 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>352</ID>
<type>DA_FROM</type>
<position>80,-101.5</position>
<input>
<ID>IN_0</ID>539 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>208</ID>
<type>DA_FROM</type>
<position>-9.5,-59.5</position>
<input>
<ID>IN_0</ID>279 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>209</ID>
<type>DA_FROM</type>
<position>-11.5,-59.5</position>
<input>
<ID>IN_0</ID>280 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>362</ID>
<type>DA_FROM</type>
<position>70.5,-91.5</position>
<input>
<ID>IN_0</ID>525 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>210</ID>
<type>DA_FROM</type>
<position>-45,-90</position>
<input>
<ID>IN_0</ID>355 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>211</ID>
<type>DA_FROM</type>
<position>-13.5,-59.5</position>
<input>
<ID>IN_0</ID>281 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>372</ID>
<type>DA_FROM</type>
<position>-45,-96</position>
<input>
<ID>IN_0</ID>356 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>212</ID>
<type>DE_TO</type>
<position>12.5,-83.5</position>
<input>
<ID>IN_0</ID>282 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec0</lparam></gate>
<gate>
<ID>213</ID>
<type>FF_GND</type>
<position>20,-66.5</position>
<output>
<ID>OUT_0</ID>283 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>366</ID>
<type>DA_FROM</type>
<position>-45,-72</position>
<input>
<ID>IN_0</ID>359 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>214</ID>
<type>DE_TO</type>
<position>-16,-73.5</position>
<input>
<ID>IN_0</ID>284 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDecOV</lparam></gate>
<gate>
<ID>215</ID>
<type>AE_FULLADDER_4BIT</type>
<position>11,-66.5</position>
<input>
<ID>IN_0</ID>274 </input>
<input>
<ID>IN_1</ID>275 </input>
<input>
<ID>IN_2</ID>276 </input>
<input>
<ID>IN_3</ID>277 </input>
<input>
<ID>IN_B_0</ID>285 </input>
<input>
<ID>IN_B_1</ID>287 </input>
<input>
<ID>IN_B_2</ID>287 </input>
<input>
<ID>IN_B_3</ID>287 </input>
<output>
<ID>OUT_0</ID>282 </output>
<output>
<ID>OUT_1</ID>288 </output>
<output>
<ID>OUT_2</ID>289 </output>
<output>
<ID>OUT_3</ID>290 </output>
<input>
<ID>carry_in</ID>283 </input>
<output>
<ID>carry_out</ID>273 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>360</ID>
<type>DA_FROM</type>
<position>-45,-94</position>
<input>
<ID>IN_0</ID>357 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>216</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-6.5,-66.5</position>
<input>
<ID>IN_0</ID>278 </input>
<input>
<ID>IN_1</ID>279 </input>
<input>
<ID>IN_2</ID>280 </input>
<input>
<ID>IN_3</ID>281 </input>
<input>
<ID>IN_B_0</ID>286 </input>
<input>
<ID>IN_B_1</ID>286 </input>
<input>
<ID>IN_B_2</ID>286 </input>
<input>
<ID>IN_B_3</ID>286 </input>
<output>
<ID>OUT_0</ID>291 </output>
<output>
<ID>OUT_1</ID>292 </output>
<output>
<ID>OUT_2</ID>293 </output>
<output>
<ID>OUT_3</ID>294 </output>
<input>
<ID>carry_in</ID>273 </input>
<output>
<ID>overflow</ID>284 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>217</ID>
<type>DA_FROM</type>
<position>8.5,-59.5</position>
<input>
<ID>IN_0</ID>275 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>370</ID>
<type>DA_FROM</type>
<position>-45,-84</position>
<input>
<ID>IN_0</ID>350 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>218</ID>
<type>DA_FROM</type>
<position>6.5,-59.5</position>
<input>
<ID>IN_0</ID>276 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>219</ID>
<type>DA_FROM</type>
<position>4.5,-59.5</position>
<input>
<ID>IN_0</ID>277 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>380</ID>
<type>DE_TO</type>
<position>-28.5,-116</position>
<input>
<ID>IN_0</ID>390 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>220</ID>
<type>EE_VDD</type>
<position>17,-60.5</position>
<output>
<ID>OUT_0</ID>285 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>221</ID>
<type>DA_FROM</type>
<position>-2.5,-59.5</position>
<input>
<ID>IN_0</ID>286 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>374</ID>
<type>AI_XOR2</type>
<position>-40,-71</position>
<input>
<ID>IN_0</ID>358 </input>
<input>
<ID>IN_1</ID>359 </input>
<output>
<ID>OUT</ID>361 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>DA_FROM</type>
<position>13,-59.5</position>
<input>
<ID>IN_0</ID>287 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>223</ID>
<type>DE_TO</type>
<position>11.5,-72.5</position>
<input>
<ID>IN_0</ID>288 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec1</lparam></gate>
<gate>
<ID>368</ID>
<type>AE_SMALL_INVERTER</type>
<position>90,-109.5</position>
<input>
<ID>IN_0</ID>528 </input>
<output>
<ID>OUT_0</ID>527 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>224</ID>
<type>DE_TO</type>
<position>10.5,-83.5</position>
<input>
<ID>IN_0</ID>289 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec2</lparam></gate>
<gate>
<ID>225</ID>
<type>DE_TO</type>
<position>9.5,-72.5</position>
<input>
<ID>IN_0</ID>290 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec3</lparam></gate>
<gate>
<ID>378</ID>
<type>AI_XOR2</type>
<position>-40,-83</position>
<input>
<ID>IN_0</ID>351 </input>
<input>
<ID>IN_1</ID>350 </input>
<output>
<ID>OUT</ID>364 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>226</ID>
<type>DE_TO</type>
<position>-5,-72.5</position>
<input>
<ID>IN_0</ID>291 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec4</lparam></gate>
<gate>
<ID>227</ID>
<type>DE_TO</type>
<position>-6,-83.5</position>
<input>
<ID>IN_0</ID>292 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec5</lparam></gate>
<gate>
<ID>260</ID>
<type>DA_FROM</type>
<position>-20.5,-108</position>
<input>
<ID>IN_0</ID>386 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>228</ID>
<type>DE_TO</type>
<position>-7,-72.5</position>
<input>
<ID>IN_0</ID>293 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec6</lparam></gate>
<gate>
<ID>229</ID>
<type>DE_TO</type>
<position>-8,-83.5</position>
<input>
<ID>IN_0</ID>294 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID IncDec7</lparam></gate>
<gate>
<ID>382</ID>
<type>AI_XOR2</type>
<position>-40,-95</position>
<input>
<ID>IN_0</ID>357 </input>
<input>
<ID>IN_1</ID>356 </input>
<output>
<ID>OUT</ID>367 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>230</ID>
<type>DA_FROM</type>
<position>39,1</position>
<input>
<ID>IN_0</ID>295 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec0</lparam></gate>
<gate>
<ID>231</ID>
<type>AA_AND2</type>
<position>-40,3</position>
<input>
<ID>IN_0</ID>297 </input>
<input>
<ID>IN_1</ID>296 </input>
<output>
<ID>OUT</ID>298 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>376</ID>
<type>AI_XOR2</type>
<position>-40,-75</position>
<input>
<ID>IN_0</ID>347 </input>
<input>
<ID>IN_1</ID>346 </input>
<output>
<ID>OUT</ID>362 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>232</ID>
<type>DA_FROM</type>
<position>-45,4</position>
<input>
<ID>IN_0</ID>297 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>233</ID>
<type>DA_FROM</type>
<position>47.5,-98.5</position>
<input>
<ID>IN_0</ID>456 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>258</ID>
<type>DA_FROM</type>
<position>28,-21</position>
<input>
<ID>IN_0</ID>408 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>234</ID>
<type>DA_FROM</type>
<position>-45,2</position>
<input>
<ID>IN_0</ID>296 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>235</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>0,-114</position>
<output>
<ID>A_equal_B</ID>373 </output>
<output>
<ID>A_greater_B</ID>371 </output>
<output>
<ID>A_less_B</ID>372 </output>
<input>
<ID>IN_0</ID>374 </input>
<input>
<ID>IN_1</ID>380 </input>
<input>
<ID>IN_2</ID>375 </input>
<input>
<ID>IN_3</ID>381 </input>
<input>
<ID>IN_B_0</ID>377 </input>
<input>
<ID>IN_B_1</ID>378 </input>
<input>
<ID>IN_B_2</ID>376 </input>
<input>
<ID>IN_B_3</ID>379 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_AND2</type>
<position>-40,-13</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>308 </input>
<output>
<ID>OUT</ID>310 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>236</ID>
<type>DE_TO</type>
<position>-35,3</position>
<input>
<ID>IN_0</ID>298 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND0</lparam></gate>
<gate>
<ID>237</ID>
<type>AA_AND2</type>
<position>-40,-1</position>
<input>
<ID>IN_0</ID>300 </input>
<input>
<ID>IN_1</ID>299 </input>
<output>
<ID>OUT</ID>301 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>262</ID>
<type>DA_FROM</type>
<position>-45,-10</position>
<input>
<ID>IN_0</ID>305 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>238</ID>
<type>DA_FROM</type>
<position>53.5,-87.5</position>
<input>
<ID>IN_0</ID>443 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>239</ID>
<type>DA_FROM</type>
<position>48.5,4.5</position>
<input>
<ID>IN_0</ID>370 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR0</lparam></gate>
<gate>
<ID>256</ID>
<type>AA_AND2</type>
<position>-40,-9</position>
<input>
<ID>IN_0</ID>306 </input>
<input>
<ID>IN_1</ID>305 </input>
<output>
<ID>OUT</ID>307 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>DA_FROM</type>
<position>-45,0</position>
<input>
<ID>IN_0</ID>300 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>241</ID>
<type>DA_FROM</type>
<position>47.5,-104.5</position>
<input>
<ID>IN_0</ID>452 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND3</lparam></gate>
<gate>
<ID>266</ID>
<type>DA_FROM</type>
<position>-3,-103</position>
<input>
<ID>IN_0</ID>380 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>242</ID>
<type>DA_FROM</type>
<position>-45,-2</position>
<input>
<ID>IN_0</ID>299 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>243</ID>
<type>DE_TO</type>
<position>-35,-1</position>
<input>
<ID>IN_0</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND1</lparam></gate>
<gate>
<ID>276</ID>
<type>AE_SMALL_INVERTER</type>
<position>42,-75</position>
<input>
<ID>IN_0</ID>425 </input>
<output>
<ID>OUT_0</ID>426 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>244</ID>
<type>DA_FROM</type>
<position>91,-69</position>
<input>
<ID>IN_0</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND6</lparam></gate>
<gate>
<ID>245</ID>
<type>AA_AND2</type>
<position>-40,-5</position>
<input>
<ID>IN_0</ID>303 </input>
<input>
<ID>IN_1</ID>302 </input>
<output>
<ID>OUT</ID>304 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>270</ID>
<type>DA_FROM</type>
<position>39,-36</position>
<input>
<ID>IN_0</ID>409 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum1</lparam></gate>
<gate>
<ID>246</ID>
<type>DA_FROM</type>
<position>81.5,-73</position>
<input>
<ID>IN_0</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum6</lparam></gate>
<gate>
<ID>247</ID>
<type>DA_FROM</type>
<position>-45,-4</position>
<input>
<ID>IN_0</ID>303 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>264</ID>
<type>DA_FROM</type>
<position>27,-56</position>
<input>
<ID>IN_0</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>248</ID>
<type>DA_FROM</type>
<position>-14.5,-103</position>
<input>
<ID>IN_0</ID>384 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>249</ID>
<type>DA_FROM</type>
<position>54.5,-15</position>
<input>
<ID>IN_0</ID>403 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>274</ID>
<type>DA_FROM</type>
<position>-45,-14</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>250</ID>
<type>DA_FROM</type>
<position>-45,-6</position>
<input>
<ID>IN_0</ID>302 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>251</ID>
<type>DE_TO</type>
<position>-35,-5</position>
<input>
<ID>IN_0</ID>304 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND2</lparam></gate>
<gate>
<ID>284</ID>
<type>DA_FROM</type>
<position>-16.5,-103</position>
<input>
<ID>IN_0</ID>385 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>252</ID>
<type>DA_FROM</type>
<position>48.5,-32</position>
<input>
<ID>IN_0</ID>412 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND1</lparam></gate>
<gate>
<ID>253</ID>
<type>DA_FROM</type>
<position>91,-98.5</position>
<input>
<ID>IN_0</ID>536 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>278</ID>
<type>DA_FROM</type>
<position>-45,-52</position>
<input>
<ID>IN_0</ID>331 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>254</ID>
<type>DA_FROM</type>
<position>-13.5,-108</position>
<input>
<ID>IN_0</ID>382 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>255</ID>
<type>AE_SMALL_INVERTER</type>
<position>43,-38</position>
<input>
<ID>IN_0</ID>405 </input>
<output>
<ID>OUT_0</ID>406 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>272</ID>
<type>DA_FROM</type>
<position>-4,-108</position>
<input>
<ID>IN_0</ID>375 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>257</ID>
<type>DA_FROM</type>
<position>96,19.5</position>
<input>
<ID>IN_0</ID>462 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>259</ID>
<type>DA_FROM</type>
<position>-45,-8</position>
<input>
<ID>IN_0</ID>306 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>261</ID>
<type>DA_FROM</type>
<position>39,-33.5</position>
<input>
<ID>IN_0</ID>411 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec1</lparam></gate>
<gate>
<ID>263</ID>
<type>DE_TO</type>
<position>-35,-9</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND3</lparam></gate>
<gate>
<ID>265</ID>
<type>DA_FROM</type>
<position>99,14.5</position>
<input>
<ID>IN_0</ID>464 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>267</ID>
<type>DA_FROM</type>
<position>27.5,-107.5</position>
<input>
<ID>IN_0</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff3</lparam></gate>
<gate>
<ID>269</ID>
<type>DA_FROM</type>
<position>82.5,-1.5</position>
<input>
<ID>IN_0</ID>469 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum4</lparam></gate>
<gate>
<ID>271</ID>
<type>DA_FROM</type>
<position>-45,-12</position>
<input>
<ID>IN_0</ID>309 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>273</ID>
<type>DA_FROM</type>
<position>36.5,-66</position>
<input>
<ID>IN_0</ID>439 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>275</ID>
<type>DE_TO</type>
<position>-35,-13</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND4</lparam></gate>
<gate>
<ID>277</ID>
<type>DA_FROM</type>
<position>91,-102.5</position>
<input>
<ID>IN_0</ID>534 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR7</lparam></gate>
<gate>
<ID>279</ID>
<type>AM_MUX_16x1</type>
<position>53,-69.5</position>
<input>
<ID>IN_0</ID>425 </input>
<input>
<ID>IN_1</ID>425 </input>
<input>
<ID>IN_10</ID>434 </input>
<input>
<ID>IN_11</ID>439 </input>
<input>
<ID>IN_12</ID>437 </input>
<input>
<ID>IN_13</ID>438 </input>
<input>
<ID>IN_14</ID>436 </input>
<input>
<ID>IN_15</ID>435 </input>
<input>
<ID>IN_2</ID>426 </input>
<input>
<ID>IN_3</ID>427 </input>
<input>
<ID>IN_4</ID>429 </input>
<input>
<ID>IN_5</ID>430 </input>
<input>
<ID>IN_6</ID>431 </input>
<input>
<ID>IN_7</ID>431 </input>
<input>
<ID>IN_8</ID>432 </input>
<input>
<ID>IN_9</ID>433 </input>
<output>
<ID>OUT</ID>420 </output>
<input>
<ID>SEL_0</ID>424 </input>
<input>
<ID>SEL_1</ID>423 </input>
<input>
<ID>SEL_2</ID>421 </input>
<input>
<ID>SEL_3</ID>422 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>281</ID>
<type>DA_FROM</type>
<position>97,-87.5</position>
<input>
<ID>IN_0</ID>523 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>283</ID>
<type>DA_FROM</type>
<position>-45,-16</position>
<input>
<ID>IN_0</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>285</ID>
<type>DA_FROM</type>
<position>51.5,-87.5</position>
<input>
<ID>IN_0</ID>442 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>287</ID>
<type>DE_TO</type>
<position>-35,-17</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND5</lparam></gate>
<gate>
<ID>289</ID>
<type>AE_SMALL_INVERTER</type>
<position>91,-2.5</position>
<input>
<ID>IN_0</ID>468 </input>
<output>
<ID>OUT_0</ID>467 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>291</ID>
<type>DA_FROM</type>
<position>71.5,13.5</position>
<input>
<ID>IN_0</ID>468 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>293</ID>
<type>DE_TO</type>
<position>102,-105</position>
<input>
<ID>IN_0</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R7</lparam></gate>
<gate>
<ID>295</ID>
<type>DA_FROM</type>
<position>-45,-20</position>
<input>
<ID>IN_0</ID>315 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>297</ID>
<type>DA_FROM</type>
<position>36.5,-68</position>
<input>
<ID>IN_0</ID>433 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR2</lparam></gate>
<gate>
<ID>299</ID>
<type>AM_MUX_16x1</type>
<position>97.5,-32.5</position>
<input>
<ID>IN_0</ID>485 </input>
<input>
<ID>IN_1</ID>485 </input>
<input>
<ID>IN_10</ID>494 </input>
<input>
<ID>IN_11</ID>499 </input>
<input>
<ID>IN_12</ID>497 </input>
<input>
<ID>IN_13</ID>498 </input>
<input>
<ID>IN_14</ID>496 </input>
<input>
<ID>IN_15</ID>495 </input>
<input>
<ID>IN_2</ID>486 </input>
<input>
<ID>IN_3</ID>487 </input>
<input>
<ID>IN_4</ID>489 </input>
<input>
<ID>IN_5</ID>490 </input>
<input>
<ID>IN_6</ID>491 </input>
<input>
<ID>IN_7</ID>491 </input>
<input>
<ID>IN_8</ID>492 </input>
<input>
<ID>IN_9</ID>493 </input>
<output>
<ID>OUT</ID>480 </output>
<input>
<ID>SEL_0</ID>484 </input>
<input>
<ID>SEL_1</ID>483 </input>
<input>
<ID>SEL_2</ID>481 </input>
<input>
<ID>SEL_3</ID>482 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>301</ID>
<type>AA_AND2</type>
<position>-40,-25</position>
<input>
<ID>IN_0</ID>318 </input>
<input>
<ID>IN_1</ID>317 </input>
<output>
<ID>OUT</ID>319 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>DA_FROM</type>
<position>92,6.5</position>
<input>
<ID>IN_0</ID>477 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>305</ID>
<type>DA_FROM</type>
<position>47.5,-67</position>
<input>
<ID>IN_0</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR2</lparam></gate>
<gate>
<ID>307</ID>
<type>DE_TO</type>
<position>-35,-25</position>
<input>
<ID>IN_0</ID>319 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND7</lparam></gate>
<gate>
<ID>309</ID>
<type>DA_FROM</type>
<position>-45,-48</position>
<input>
<ID>IN_0</ID>328 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>311</ID>
<type>DA_FROM</type>
<position>-45,-32</position>
<input>
<ID>IN_0</ID>321 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>313</ID>
<type>DA_FROM</type>
<position>71.5,-21</position>
<input>
<ID>IN_0</ID>488 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>315</ID>
<type>DA_FROM</type>
<position>-45,-38</position>
<input>
<ID>IN_0</ID>323 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>317</ID>
<type>DA_FROM</type>
<position>-45,-56</position>
<input>
<ID>IN_0</ID>332 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>319</ID>
<type>AE_OR2</type>
<position>-40,-41</position>
<input>
<ID>IN_0</ID>325 </input>
<input>
<ID>IN_1</ID>324 </input>
<output>
<ID>OUT</ID>338 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>320</ID>
<type>DA_FROM</type>
<position>-45,-42</position>
<input>
<ID>IN_0</ID>324 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>321</ID>
<type>DA_FROM</type>
<position>-45,-44</position>
<input>
<ID>IN_0</ID>326 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>322</ID>
<type>AE_OR2</type>
<position>-40,-57</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>333 </input>
<output>
<ID>OUT</ID>342 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>323</ID>
<type>DA_FROM</type>
<position>-45,-46</position>
<input>
<ID>IN_0</ID>327 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>324</ID>
<type>DA_FROM</type>
<position>80,-66</position>
<input>
<ID>IN_0</ID>519 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>325</ID>
<type>DA_FROM</type>
<position>-45,-50</position>
<input>
<ID>IN_0</ID>329 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y4</lparam></gate>
<gate>
<ID>326</ID>
<type>AM_MUX_16x1</type>
<position>96.5,-69.5</position>
<input>
<ID>IN_0</ID>505 </input>
<input>
<ID>IN_1</ID>505 </input>
<input>
<ID>IN_10</ID>514 </input>
<input>
<ID>IN_11</ID>519 </input>
<input>
<ID>IN_12</ID>517 </input>
<input>
<ID>IN_13</ID>518 </input>
<input>
<ID>IN_14</ID>516 </input>
<input>
<ID>IN_15</ID>515 </input>
<input>
<ID>IN_2</ID>506 </input>
<input>
<ID>IN_3</ID>507 </input>
<input>
<ID>IN_4</ID>509 </input>
<input>
<ID>IN_5</ID>510 </input>
<input>
<ID>IN_6</ID>511 </input>
<input>
<ID>IN_7</ID>511 </input>
<input>
<ID>IN_8</ID>512 </input>
<input>
<ID>IN_9</ID>513 </input>
<output>
<ID>OUT</ID>500 </output>
<input>
<ID>SEL_0</ID>504 </input>
<input>
<ID>SEL_1</ID>503 </input>
<input>
<ID>SEL_2</ID>501 </input>
<input>
<ID>SEL_3</ID>502 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>327</ID>
<type>DA_FROM</type>
<position>-45,-54</position>
<input>
<ID>IN_0</ID>330 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y5</lparam></gate>
<gate>
<ID>328</ID>
<type>DA_FROM</type>
<position>95,-87.5</position>
<input>
<ID>IN_0</ID>522 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>329</ID>
<type>DA_FROM</type>
<position>-45,-58</position>
<input>
<ID>IN_0</ID>333 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>330</ID>
<type>DA_FROM</type>
<position>71,-72</position>
<input>
<ID>IN_0</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff6</lparam></gate>
<gate>
<ID>331</ID>
<type>DA_FROM</type>
<position>-45,-62</position>
<input>
<ID>IN_0</ID>335 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>332</ID>
<type>DA_FROM</type>
<position>72,-35</position>
<input>
<ID>IN_0</ID>490 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff5</lparam></gate>
<gate>
<ID>333</ID>
<type>AE_OR2</type>
<position>-40,-33</position>
<input>
<ID>IN_0</ID>321 </input>
<input>
<ID>IN_1</ID>320 </input>
<output>
<ID>OUT</ID>336 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>334</ID>
<type>DA_FROM</type>
<position>91,-63</position>
<input>
<ID>IN_0</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>335</ID>
<type>DA_FROM</type>
<position>80,-97.5</position>
<input>
<ID>IN_0</ID>535 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>336</ID>
<type>AE_OR2</type>
<position>-40,-37</position>
<input>
<ID>IN_0</ID>322 </input>
<input>
<ID>IN_1</ID>323 </input>
<output>
<ID>OUT</ID>337 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>337</ID>
<type>AE_OR2</type>
<position>-40,-45</position>
<input>
<ID>IN_0</ID>326 </input>
<input>
<ID>IN_1</ID>327 </input>
<output>
<ID>OUT</ID>339 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>338</ID>
<type>DA_FROM</type>
<position>92,-28</position>
<input>
<ID>IN_0</ID>497 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>339</ID>
<type>AE_OR2</type>
<position>-40,-49</position>
<input>
<ID>IN_0</ID>328 </input>
<input>
<ID>IN_1</ID>329 </input>
<output>
<ID>OUT</ID>340 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>340</ID>
<type>DA_FROM</type>
<position>98,-92.5</position>
<input>
<ID>IN_0</ID>524 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>341</ID>
<type>DA_FROM</type>
<position>70.5,-93.5</position>
<input>
<ID>IN_0</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y7</lparam></gate>
<gate>
<ID>342</ID>
<type>AE_OR2</type>
<position>-40,-53</position>
<input>
<ID>IN_0</ID>331 </input>
<input>
<ID>IN_1</ID>330 </input>
<output>
<ID>OUT</ID>341 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>343</ID>
<type>AE_OR2</type>
<position>-40,-61</position>
<input>
<ID>IN_0</ID>334 </input>
<input>
<ID>IN_1</ID>335 </input>
<output>
<ID>OUT</ID>343 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>345</ID>
<type>DA_FROM</type>
<position>81.5,-108.5</position>
<input>
<ID>IN_0</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum7</lparam></gate>
<gate>
<ID>347</ID>
<type>DA_FROM</type>
<position>80,-68</position>
<input>
<ID>IN_0</ID>513 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR6</lparam></gate>
<gate>
<ID>348</ID>
<type>DE_TO</type>
<position>-35,-37</position>
<input>
<ID>IN_0</ID>337 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR1</lparam></gate>
<gate>
<ID>349</ID>
<type>DE_TO</type>
<position>-35,-41</position>
<input>
<ID>IN_0</ID>338 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR2</lparam></gate>
<gate>
<ID>351</ID>
<type>DE_TO</type>
<position>-35,-45</position>
<input>
<ID>IN_0</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR3</lparam></gate>
<gate>
<ID>353</ID>
<type>DA_FROM</type>
<position>81,-27</position>
<input>
<ID>IN_0</ID>498 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>355</ID>
<type>DE_TO</type>
<position>-35,-57</position>
<input>
<ID>IN_0</ID>342 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR6</lparam></gate>
<gate>
<ID>357</ID>
<type>DE_TO</type>
<position>-35,-61</position>
<input>
<ID>IN_0</ID>343 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR7</lparam></gate>
<gate>
<ID>359</ID>
<type>DA_FROM</type>
<position>91,-100.5</position>
<input>
<ID>IN_0</ID>537 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>361</ID>
<type>DA_FROM</type>
<position>-45,-82</position>
<input>
<ID>IN_0</ID>351 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>363</ID>
<type>DA_FROM</type>
<position>-45,-66</position>
<input>
<ID>IN_0</ID>344 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>365</ID>
<type>AE_SMALL_INVERTER</type>
<position>85.5,-75</position>
<input>
<ID>IN_0</ID>505 </input>
<output>
<ID>OUT_0</ID>506 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>367</ID>
<type>DA_FROM</type>
<position>-45,-74</position>
<input>
<ID>IN_0</ID>347 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>369</ID>
<type>DA_FROM</type>
<position>-45,-78</position>
<input>
<ID>IN_0</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>371</ID>
<type>DA_FROM</type>
<position>-45,-92</position>
<input>
<ID>IN_0</ID>354 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>373</ID>
<type>AI_XOR2</type>
<position>-40,-67</position>
<input>
<ID>IN_0</ID>344 </input>
<input>
<ID>IN_1</ID>345 </input>
<output>
<ID>OUT</ID>360 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>375</ID>
<type>DA_FROM</type>
<position>96,-92.5</position>
<input>
<ID>IN_0</ID>521 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>377</ID>
<type>AI_XOR2</type>
<position>-40,-79</position>
<input>
<ID>IN_0</ID>348 </input>
<input>
<ID>IN_1</ID>349 </input>
<output>
<ID>OUT</ID>363 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>379</ID>
<type>AI_XOR2</type>
<position>-40,-87</position>
<input>
<ID>IN_0</ID>353 </input>
<input>
<ID>IN_1</ID>352 </input>
<output>
<ID>OUT</ID>365 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>381</ID>
<type>AI_XOR2</type>
<position>-40,-91</position>
<input>
<ID>IN_0</ID>355 </input>
<input>
<ID>IN_1</ID>354 </input>
<output>
<ID>OUT</ID>366 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>383</ID>
<type>DE_TO</type>
<position>-35,-67</position>
<input>
<ID>IN_0</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR0</lparam></gate>
<gate>
<ID>384</ID>
<type>DE_TO</type>
<position>-35,-71</position>
<input>
<ID>IN_0</ID>361 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR1</lparam></gate>
<gate>
<ID>385</ID>
<type>DE_TO</type>
<position>-35,-75</position>
<input>
<ID>IN_0</ID>362 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR2</lparam></gate>
<gate>
<ID>386</ID>
<type>DE_TO</type>
<position>-35,-79</position>
<input>
<ID>IN_0</ID>363 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR3</lparam></gate>
<gate>
<ID>387</ID>
<type>DA_FROM</type>
<position>81.5,-70.5</position>
<input>
<ID>IN_0</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec6</lparam></gate>
<gate>
<ID>388</ID>
<type>DE_TO</type>
<position>-35,-83</position>
<input>
<ID>IN_0</ID>364 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR4</lparam></gate>
<gate>
<ID>389</ID>
<type>DA_FROM</type>
<position>36.5,-64</position>
<input>
<ID>IN_0</ID>438 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>390</ID>
<type>DA_FROM</type>
<position>48.5,6.5</position>
<input>
<ID>IN_0</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>391</ID>
<type>DE_TO</type>
<position>-35,-87</position>
<input>
<ID>IN_0</ID>365 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR5</lparam></gate>
<gate>
<ID>392</ID>
<type>DE_TO</type>
<position>-35,-91</position>
<input>
<ID>IN_0</ID>366 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR6</lparam></gate>
<gate>
<ID>393</ID>
<type>AE_OR2</type>
<position>-39.5,-112</position>
<input>
<ID>IN_0</ID>391 </input>
<input>
<ID>IN_1</ID>392 </input>
<output>
<ID>OUT</ID>393 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>394</ID>
<type>DE_TO</type>
<position>-35,-95</position>
<input>
<ID>IN_0</ID>367 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR7</lparam></gate>
<gate>
<ID>395</ID>
<type>DE_TO</type>
<position>58.5,-105</position>
<input>
<ID>IN_0</ID>440 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R3</lparam></gate>
<gate>
<ID>396</ID>
<type>DA_FROM</type>
<position>-15.5,-108</position>
<input>
<ID>IN_0</ID>383 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y6</lparam></gate>
<gate>
<ID>397</ID>
<type>DA_FROM</type>
<position>48.5,2.5</position>
<input>
<ID>IN_0</ID>368 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND0</lparam></gate>
<gate>
<ID>398</ID>
<type>DA_FROM</type>
<position>37.5,3.5</position>
<input>
<ID>IN_0</ID>369 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR0</lparam></gate>
<gate>
<ID>399</ID>
<type>DE_TO</type>
<position>-44.5,-116</position>
<input>
<ID>IN_0</ID>394 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>400</ID>
<type>DA_FROM</type>
<position>47.5,-102.5</position>
<input>
<ID>IN_0</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR3</lparam></gate>
<gate>
<ID>401</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>-18.5,-114</position>
<output>
<ID>A_equal_B</ID>391 </output>
<output>
<ID>A_greater_B</ID>392 </output>
<output>
<ID>A_less_B</ID>390 </output>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>389 </input>
<input>
<ID>IN_2</ID>387 </input>
<input>
<ID>IN_3</ID>388 </input>
<input>
<ID>IN_B_0</ID>382 </input>
<input>
<ID>IN_B_1</ID>384 </input>
<input>
<ID>IN_B_2</ID>383 </input>
<input>
<ID>IN_B_3</ID>385 </input>
<input>
<ID>in_A_equal_B</ID>373 </input>
<input>
<ID>in_A_greater_B</ID>371 </input>
<input>
<ID>in_A_less_B</ID>372 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>402</ID>
<type>DA_FROM</type>
<position>37.5,5.5</position>
<input>
<ID>IN_0</ID>399 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>403</ID>
<type>DA_FROM</type>
<position>2,-103</position>
<input>
<ID>IN_0</ID>379 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>404</ID>
<type>DA_FROM</type>
<position>98,-15</position>
<input>
<ID>IN_0</ID>483 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>405</ID>
<type>DA_FROM</type>
<position>48.5,8.5</position>
<input>
<ID>IN_0</ID>396 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>406</ID>
<type>DA_FROM</type>
<position>3,-108</position>
<input>
<ID>IN_0</ID>376 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>407</ID>
<type>DA_FROM</type>
<position>-22.5,-108</position>
<input>
<ID>IN_0</ID>387 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X6</lparam></gate>
<gate>
<ID>408</ID>
<type>DA_FROM</type>
<position>92,4.5</position>
<input>
<ID>IN_0</ID>474 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR4</lparam></gate>
<gate>
<ID>409</ID>
<type>DA_FROM</type>
<position>98,-57</position>
<input>
<ID>IN_0</ID>504 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>410</ID>
<type>DA_FROM</type>
<position>-21.5,-103</position>
<input>
<ID>IN_0</ID>389 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>411</ID>
<type>DA_FROM</type>
<position>37.5,9.5</position>
<input>
<ID>IN_0</ID>395 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>412</ID>
<type>AE_SMALL_INVERTER</type>
<position>86.5,-38</position>
<input>
<ID>IN_0</ID>485 </input>
<output>
<ID>OUT_0</ID>486 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>413</ID>
<type>DA_FROM</type>
<position>-23.5,-103</position>
<input>
<ID>IN_0</ID>388 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X7</lparam></gate>
<gate>
<ID>414</ID>
<type>DA_FROM</type>
<position>52.5,-15</position>
<input>
<ID>IN_0</ID>402 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>415</ID>
<type>DA_FROM</type>
<position>-2,-108</position>
<input>
<ID>IN_0</ID>374 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>416</ID>
<type>DA_FROM</type>
<position>82.5,-33.5</position>
<input>
<ID>IN_0</ID>491 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec5</lparam></gate>
<gate>
<ID>417</ID>
<type>DE_TO</type>
<position>59.5,-32.5</position>
<input>
<ID>IN_0</ID>400 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1</lparam></gate>
<gate>
<ID>418</ID>
<type>DA_FROM</type>
<position>4,-103</position>
<input>
<ID>IN_0</ID>378 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>419</ID>
<type>DA_FROM</type>
<position>-5,-103</position>
<input>
<ID>IN_0</ID>381 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>420</ID>
<type>DA_FROM</type>
<position>37.5,7.5</position>
<input>
<ID>IN_0</ID>398 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>421</ID>
<type>DA_FROM</type>
<position>71,-107.5</position>
<input>
<ID>IN_0</ID>530 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff7</lparam></gate>
<gate>
<ID>422</ID>
<type>DE_TO</type>
<position>-28.5,-112</position>
<input>
<ID>IN_0</ID>392 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>423</ID>
<type>DE_TO</type>
<position>-31.5,-114</position>
<input>
<ID>IN_0</ID>391 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>424</ID>
<type>DA_FROM</type>
<position>96,-57</position>
<input>
<ID>IN_0</ID>501 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>425</ID>
<type>AE_OR2</type>
<position>-39.5,-116</position>
<input>
<ID>IN_0</ID>390 </input>
<input>
<ID>IN_1</ID>391 </input>
<output>
<ID>OUT</ID>394 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>426</ID>
<type>DE_TO</type>
<position>-44.5,-112</position>
<input>
<ID>IN_0</ID>393 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>427</ID>
<type>DA_FROM</type>
<position>98,19.5</position>
<input>
<ID>IN_0</ID>463 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>428</ID>
<type>DA_FROM</type>
<position>97,-20</position>
<input>
<ID>IN_0</ID>481 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>429</ID>
<type>DA_FROM</type>
<position>92,8.5</position>
<input>
<ID>IN_0</ID>476 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>430</ID>
<type>AE_SMALL_INVERTER</type>
<position>91,-37</position>
<input>
<ID>IN_0</ID>488 </input>
<output>
<ID>OUT_0</ID>487 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>431</ID>
<type>DA_FROM</type>
<position>72,-0.5</position>
<input>
<ID>IN_0</ID>470 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff4</lparam></gate>
<gate>
<ID>432</ID>
<type>DA_FROM</type>
<position>28,-19</position>
<input>
<ID>IN_0</ID>405 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>433</ID>
<type>AM_MUX_16x1</type>
<position>54,-32.5</position>
<input>
<ID>IN_0</ID>405 </input>
<input>
<ID>IN_1</ID>405 </input>
<input>
<ID>IN_10</ID>414 </input>
<input>
<ID>IN_11</ID>419 </input>
<input>
<ID>IN_12</ID>417 </input>
<input>
<ID>IN_13</ID>418 </input>
<input>
<ID>IN_14</ID>416 </input>
<input>
<ID>IN_15</ID>415 </input>
<input>
<ID>IN_2</ID>406 </input>
<input>
<ID>IN_3</ID>407 </input>
<input>
<ID>IN_4</ID>409 </input>
<input>
<ID>IN_5</ID>410 </input>
<input>
<ID>IN_6</ID>411 </input>
<input>
<ID>IN_7</ID>411 </input>
<input>
<ID>IN_8</ID>412 </input>
<input>
<ID>IN_9</ID>413 </input>
<output>
<ID>OUT</ID>400 </output>
<input>
<ID>SEL_0</ID>404 </input>
<input>
<ID>SEL_1</ID>403 </input>
<input>
<ID>SEL_2</ID>401 </input>
<input>
<ID>SEL_3</ID>402 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>434</ID>
<type>DA_FROM</type>
<position>55.5,-20</position>
<input>
<ID>IN_0</ID>404 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>435</ID>
<type>DA_FROM</type>
<position>53.5,-20</position>
<input>
<ID>IN_0</ID>401 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>436</ID>
<type>DA_FROM</type>
<position>27,-93.5</position>
<input>
<ID>IN_0</ID>448 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>437</ID>
<type>AE_SMALL_INVERTER</type>
<position>47.5,-37</position>
<input>
<ID>IN_0</ID>408 </input>
<output>
<ID>OUT_0</ID>407 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>438</ID>
<type>DA_FROM</type>
<position>28.5,-35</position>
<input>
<ID>IN_0</ID>410 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff1</lparam></gate>
<gate>
<ID>439</ID>
<type>DA_FROM</type>
<position>48.5,-30</position>
<input>
<ID>IN_0</ID>414 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR1</lparam></gate>
<gate>
<ID>440</ID>
<type>DA_FROM</type>
<position>37.5,-31</position>
<input>
<ID>IN_0</ID>413 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR1</lparam></gate>
<gate>
<ID>441</ID>
<type>DA_FROM</type>
<position>48.5,-28</position>
<input>
<ID>IN_0</ID>417 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>442</ID>
<type>DA_FROM</type>
<position>37.5,-27</position>
<input>
<ID>IN_0</ID>418 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>443</ID>
<type>DA_FROM</type>
<position>37.5,-29</position>
<input>
<ID>IN_0</ID>419 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>444</ID>
<type>DE_TO</type>
<position>58.5,-69.5</position>
<input>
<ID>IN_0</ID>420 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R2</lparam></gate>
<gate>
<ID>445</ID>
<type>DA_FROM</type>
<position>36.5,-97.5</position>
<input>
<ID>IN_0</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>446</ID>
<type>DA_FROM</type>
<position>53.5,-52</position>
<input>
<ID>IN_0</ID>423 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>447</ID>
<type>DA_FROM</type>
<position>51.5,-52</position>
<input>
<ID>IN_0</ID>422 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>448</ID>
<type>AE_SMALL_INVERTER</type>
<position>46.5,-74</position>
<input>
<ID>IN_0</ID>428 </input>
<output>
<ID>OUT_0</ID>427 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>449</ID>
<type>DA_FROM</type>
<position>27.5,-72</position>
<input>
<ID>IN_0</ID>430 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Diff2</lparam></gate>
<gate>
<ID>450</ID>
<type>DA_FROM</type>
<position>36.5,-103.5</position>
<input>
<ID>IN_0</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR3</lparam></gate>
<gate>
<ID>451</ID>
<type>DA_FROM</type>
<position>47.5,-63</position>
<input>
<ID>IN_0</ID>436 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>452</ID>
<type>DA_FROM</type>
<position>27,-91.5</position>
<input>
<ID>IN_0</ID>445 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>453</ID>
<type>DA_FROM</type>
<position>54.5,-92.5</position>
<input>
<ID>IN_0</ID>444 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>454</ID>
<type>DA_FROM</type>
<position>52.5,-92.5</position>
<input>
<ID>IN_0</ID>441 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>455</ID>
<type>AE_SMALL_INVERTER</type>
<position>42,-110.5</position>
<input>
<ID>IN_0</ID>445 </input>
<output>
<ID>OUT_0</ID>446 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>456</ID>
<type>AE_SMALL_INVERTER</type>
<position>46.5,-109.5</position>
<input>
<ID>IN_0</ID>448 </input>
<output>
<ID>OUT_0</ID>447 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>457</ID>
<type>DA_FROM</type>
<position>38,-108.5</position>
<input>
<ID>IN_0</ID>449 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum3</lparam></gate>
<gate>
<ID>458</ID>
<type>DA_FROM</type>
<position>38,-106</position>
<input>
<ID>IN_0</ID>451 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec3</lparam></gate>
<gate>
<ID>459</ID>
<type>DA_FROM</type>
<position>47.5,-100.5</position>
<input>
<ID>IN_0</ID>457 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>460</ID>
<type>DA_FROM</type>
<position>36.5,-99.5</position>
<input>
<ID>IN_0</ID>458 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>461</ID>
<type>DA_FROM</type>
<position>36.5,-101.5</position>
<input>
<ID>IN_0</ID>459 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>462</ID>
<type>DA_FROM</type>
<position>71.5,15.5</position>
<input>
<ID>IN_0</ID>465 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X4</lparam></gate>
<gate>
<ID>463</ID>
<type>DE_TO</type>
<position>103,2</position>
<input>
<ID>IN_0</ID>460 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R4</lparam></gate>
<gate>
<ID>464</ID>
<type>DA_FROM</type>
<position>81,-25</position>
<input>
<ID>IN_0</ID>495 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>465</ID>
<type>AM_MUX_16x1</type>
<position>97.5,2</position>
<input>
<ID>IN_0</ID>465 </input>
<input>
<ID>IN_1</ID>465 </input>
<input>
<ID>IN_10</ID>474 </input>
<input>
<ID>IN_11</ID>479 </input>
<input>
<ID>IN_12</ID>477 </input>
<input>
<ID>IN_13</ID>478 </input>
<input>
<ID>IN_14</ID>476 </input>
<input>
<ID>IN_15</ID>475 </input>
<input>
<ID>IN_2</ID>466 </input>
<input>
<ID>IN_3</ID>467 </input>
<input>
<ID>IN_4</ID>469 </input>
<input>
<ID>IN_5</ID>470 </input>
<input>
<ID>IN_6</ID>471 </input>
<input>
<ID>IN_7</ID>471 </input>
<input>
<ID>IN_8</ID>472 </input>
<input>
<ID>IN_9</ID>473 </input>
<output>
<ID>OUT</ID>460 </output>
<input>
<ID>SEL_0</ID>464 </input>
<input>
<ID>SEL_1</ID>463 </input>
<input>
<ID>SEL_2</ID>461 </input>
<input>
<ID>SEL_3</ID>462 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>466</ID>
<type>DA_FROM</type>
<position>91,-65</position>
<input>
<ID>IN_0</ID>517 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ></lparam></gate>
<gate>
<ID>467</ID>
<type>DA_FROM</type>
<position>97,14.5</position>
<input>
<ID>IN_0</ID>461 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>468</ID>
<type>AE_SMALL_INVERTER</type>
<position>86.5,-3.5</position>
<input>
<ID>IN_0</ID>465 </input>
<output>
<ID>OUT_0</ID>466 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>469</ID>
<type>DA_FROM</type>
<position>82.5,1</position>
<input>
<ID>IN_0</ID>471 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec4</lparam></gate>
<gate>
<ID>470</ID>
<type>DA_FROM</type>
<position>91,-104.5</position>
<input>
<ID>IN_0</ID>532 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND7</lparam></gate>
<gate>
<ID>471</ID>
<type>DA_FROM</type>
<position>92,2.5</position>
<input>
<ID>IN_0</ID>472 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND4</lparam></gate>
<gate>
<ID>472</ID>
<type>DA_FROM</type>
<position>81,3.5</position>
<input>
<ID>IN_0</ID>473 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR4</lparam></gate>
<gate>
<ID>473</ID>
<type>DA_FROM</type>
<position>81,7.5</position>
<input>
<ID>IN_0</ID>478 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>474</ID>
<type>DA_FROM</type>
<position>71.5,-19</position>
<input>
<ID>IN_0</ID>485 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X5</lparam></gate>
<gate>
<ID>476</ID>
<type>DA_FROM</type>
<position>99,-20</position>
<input>
<ID>IN_0</ID>484 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C0</lparam></gate>
<gate>
<ID>477</ID>
<type>DA_FROM</type>
<position>96,-15</position>
<input>
<ID>IN_0</ID>482 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>478</ID>
<type>DA_FROM</type>
<position>82.5,-36</position>
<input>
<ID>IN_0</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum5</lparam></gate>
<gate>
<ID>479</ID>
<type>DA_FROM</type>
<position>92,-30</position>
<input>
<ID>IN_0</ID>494 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID XOR5</lparam></gate>
<gate>
<ID>480</ID>
<type>DA_FROM</type>
<position>92,-32</position>
<input>
<ID>IN_0</ID>492 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND5</lparam></gate>
<gate>
<ID>482</ID>
<type>DA_FROM</type>
<position>92,-26</position>
<input>
<ID>IN_0</ID>496 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID </lparam></gate>
<gate>
<ID>483</ID>
<type>DA_FROM</type>
<position>81,-29</position>
<input>
<ID>IN_0</ID>499 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID >=</lparam></gate>
<gate>
<ID>484</ID>
<type>DE_TO</type>
<position>102,-69.5</position>
<input>
<ID>IN_0</ID>500 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R6</lparam></gate>
<gate>
<ID>486</ID>
<type>DA_FROM</type>
<position>95,-52</position>
<input>
<ID>IN_0</ID>502 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>487</ID>
<type>AE_SMALL_INVERTER</type>
<position>90,-74</position>
<input>
<ID>IN_0</ID>508 </input>
<output>
<ID>OUT_0</ID>507 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>488</ID>
<type>DA_FROM</type>
<position>80,-103.5</position>
<input>
<ID>IN_0</ID>533 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR7</lparam></gate>
<gate>
<ID>489</ID>
<type>DA_FROM</type>
<position>80,-62</position>
<input>
<ID>IN_0</ID>515 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>490</ID>
<type>AM_MUX_16x1</type>
<position>96.5,-105</position>
<input>
<ID>IN_0</ID>525 </input>
<input>
<ID>IN_1</ID>525 </input>
<input>
<ID>IN_10</ID>534 </input>
<input>
<ID>IN_11</ID>539 </input>
<input>
<ID>IN_12</ID>537 </input>
<input>
<ID>IN_13</ID>538 </input>
<input>
<ID>IN_14</ID>536 </input>
<input>
<ID>IN_15</ID>535 </input>
<input>
<ID>IN_2</ID>526 </input>
<input>
<ID>IN_3</ID>527 </input>
<input>
<ID>IN_4</ID>529 </input>
<input>
<ID>IN_5</ID>530 </input>
<input>
<ID>IN_6</ID>531 </input>
<input>
<ID>IN_7</ID>531 </input>
<input>
<ID>IN_8</ID>532 </input>
<input>
<ID>IN_9</ID>533 </input>
<output>
<ID>OUT</ID>520 </output>
<input>
<ID>SEL_0</ID>524 </input>
<input>
<ID>SEL_1</ID>523 </input>
<input>
<ID>SEL_2</ID>521 </input>
<input>
<ID>SEL_3</ID>522 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>491</ID>
<type>AE_SMALL_INVERTER</type>
<position>85.5,-110.5</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>492</ID>
<type>DA_FROM</type>
<position>81.5,-106</position>
<input>
<ID>IN_0</ID>531 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IncDec7</lparam></gate>
<gate>
<ID>493</ID>
<type>DA_FROM</type>
<position>80,-99.5</position>
<input>
<ID>IN_0</ID>538 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<wire>
<ID>416 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-26,51,-26</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>480 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>100.5,-32.5,101,-32.5</points>
<connection>
<GID>299</GID>
<name>OUT</name></connection>
<connection>
<GID>475</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>223 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-8,8,-7.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>9.5,-7.5,9.5,-7</points>
<connection>
<GID>189</GID>
<name>OUT_3</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>8,-7.5,9.5,-7.5</points>
<intersection>8 0</intersection>
<intersection>9.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>368 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>50.5,2.5,51,2.5</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>432 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-69,50,-69</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>415 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-25,51,-25</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>459 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-101.5,50,-101.5</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>395 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,9.5,51,9.5</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>267 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-5.5,40,15.5</points>
<intersection>-5.5 1</intersection>
<intersection>-4.5 4</intersection>
<intersection>-3.5 6</intersection>
<intersection>15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-5.5,51,-5.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,15.5,40,15.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>40,-4.5,51,-4.5</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>40,-3.5,41,-3.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>259 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,-27,-3.5,-25.5</points>
<connection>
<GID>186</GID>
<name>IN_1</name></connection>
<intersection>-25.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-3.5,-25.5,-2.5,-25.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>334 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-60,-43,-60</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<connection>
<GID>343</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>398 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,7.5,51,7.5</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>245 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-40.5,-5.5,-40</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>-40 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-6,-40,-6,-39.5</points>
<connection>
<GID>174</GID>
<name>OUT_1</name></connection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-6,-40,-5.5,-40</points>
<intersection>-6 1</intersection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>270 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-2.5,41.5,13.5</points>
<intersection>-2.5 1</intersection>
<intersection>13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-2.5,45.5,-2.5</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,13.5,41.5,13.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>429 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-73,50,-73</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>198 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>57,2,57.5,2</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<connection>
<GID>127</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>493 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-31,94.5,-31</points>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<connection>
<GID>299</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>233 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-31.5,8,-31</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>8.5,-31,8.5,-30.5</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>8,-31,8.5,-31</points>
<intersection>8 0</intersection>
<intersection>8.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>258 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-27,-4.5,-25.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>534 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>93,-102.5,93.5,-102.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>204 </ID>
<shape>
<vsegment>
<ID>1</ID>
<points>19.5,1,19.5,2</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>16,1,19.5,1</points>
<connection>
<GID>189</GID>
<name>IN_B_0</name></connection>
<intersection>19.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>316 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-21,-37,-21</points>
<connection>
<GID>292</GID>
<name>OUT</name></connection>
<connection>
<GID>298</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>508 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-74,84,-58</points>
<intersection>-74 1</intersection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-74,88,-74</points>
<connection>
<GID>487</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72.5,-58,84,-58</points>
<connection>
<GID>485</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>421 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-60,52.5,-59</points>
<connection>
<GID>279</GID>
<name>SEL_2</name></connection>
<connection>
<GID>126</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>261 </ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-0.5,-26.5,-0.5,-25.5</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-2.5,-26.5,-0.5,-26.5</points>
<intersection>-2.5 3</intersection>
<intersection>-0.5 1</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2.5,-27,-2.5,-26.5</points>
<connection>
<GID>186</GID>
<name>IN_2</name></connection>
<intersection>-26.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>370 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>50.5,4.5,51,4.5</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>217 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,1,-9.5,2</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<connection>
<GID>146</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>271 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-1.5,51,-1.5</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>399 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,5.5,51,5.5</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>269 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-2.5,51,-2.5</points>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>397 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>50.5,6.5,51,6.5</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>235 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-31,4.5,-30.5</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>6,-31.5,6,-31</points>
<connection>
<GID>173</GID>
<name>IN_3</name></connection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-31,6,-31</points>
<intersection>4.5 0</intersection>
<intersection>6 1</intersection></hsegment></shape></wire>
<wire>
<ID>268 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-3.5,51,-3.5</points>
<connection>
<GID>198</GID>
<name>OUT_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>396 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>50.5,8.5,51,8.5</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>255 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-27,14,-25.5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>-25.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>14,-25.5,15,-25.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>272 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-0.5,51,-0.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>248 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-41,-14.5,-36.5</points>
<connection>
<GID>174</GID>
<name>overflow</name></connection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-14.5,-41,-13,-41</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>295 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,1,51,1</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>51 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>51,0.5,51,1.5</points>
<connection>
<GID>130</GID>
<name>IN_7</name></connection>
<connection>
<GID>130</GID>
<name>IN_6</name></connection>
<intersection>1 1</intersection></vsegment></shape></wire>
<wire>
<ID>202 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>55.5,11.5,55.5,12.5</points>
<connection>
<GID>130</GID>
<name>SEL_0</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>369 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,3.5,51,3.5</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>354 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-92,-43,-92</points>
<connection>
<GID>371</GID>
<name>IN_0</name></connection>
<connection>
<GID>381</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>201 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,11.5,54.5,17.5</points>
<connection>
<GID>130</GID>
<name>SEL_1</name></connection>
<connection>
<GID>136</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>521 </ID>
<shape>
<vsegment>
<ID>4</ID>
<points>96,-95.5,96,-94.5</points>
<connection>
<GID>490</GID>
<name>SEL_2</name></connection>
<connection>
<GID>375</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>344 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-66,-43,-66</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<connection>
<GID>373</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>199 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>53.5,11.5,53.5,12.5</points>
<connection>
<GID>130</GID>
<name>SEL_2</name></connection>
<connection>
<GID>137</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>311 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-18,-43,-18</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<connection>
<GID>280</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>530 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-107.5,93.5,-107.5</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>200 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,11.5,52.5,17.5</points>
<connection>
<GID>130</GID>
<name>SEL_3</name></connection>
<connection>
<GID>139</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>315 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-20,-43,-20</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<connection>
<GID>295</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>314 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-22,-43,-22</points>
<connection>
<GID>292</GID>
<name>IN_1</name></connection>
<connection>
<GID>296</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>437 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-65,50,-65</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>206 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,1,14,2</points>
<connection>
<GID>189</GID>
<name>IN_B_2</name></connection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>14,2,15.5,2</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>447 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-109.5,50,-109.5</points>
<connection>
<GID>456</GID>
<name>OUT_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>538 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-99.5,93.5,-99.5</points>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>208 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,1,9,1.5</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>1.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>10.5,1.5,10.5,2</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>9,1.5,10.5,1.5</points>
<intersection>9 0</intersection>
<intersection>10.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>312 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-16,-43,-16</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<connection>
<GID>283</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>377 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-110,5,-110</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<connection>
<GID>235</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>520 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99.5,-105,100,-105</points>
<connection>
<GID>490</GID>
<name>OUT</name></connection>
<connection>
<GID>293</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>313 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-17,-37,-17</points>
<connection>
<GID>280</GID>
<name>OUT</name></connection>
<connection>
<GID>287</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>360 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-67,-37,-67</points>
<connection>
<GID>373</GID>
<name>OUT</name></connection>
<connection>
<GID>383</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>537 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93,-100.5,93.5,-100.5</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>215 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,1,-4.5,2</points>
<connection>
<GID>190</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>143</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>424 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-60,54.5,-59</points>
<connection>
<GID>279</GID>
<name>SEL_0</name></connection>
<connection>
<GID>138</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>256 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>16,-27,19,-27</points>
<connection>
<GID>183</GID>
<name>IN_3</name></connection>
<intersection>19 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19,-27,19,-25.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>-27 2</intersection></vsegment></shape></wire>
<wire>
<ID>239 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-31.5,-13.5,-30.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-13.5,-31.5,-11.5,-31.5</points>
<connection>
<GID>174</GID>
<name>IN_3</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>428 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-74,40.5,-58</points>
<intersection>-74 1</intersection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-74,44.5,-74</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-58,40.5,-58</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>445 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-112.5,39,-91.5</points>
<intersection>-112.5 1</intersection>
<intersection>-111.5 4</intersection>
<intersection>-110.5 7</intersection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-112.5,50,-112.5</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-91.5,39,-91.5</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>39,-111.5,50,-111.5</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>39,-110.5,40,-110.5</points>
<connection>
<GID>455</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>214 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,1,-3.5,2</points>
<connection>
<GID>190</GID>
<name>IN_B_2</name></connection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-3.5,2,-2.5,2</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>431 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-70.5,50,-70.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>50 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50,-71,50,-70</points>
<connection>
<GID>279</GID>
<name>IN_7</name></connection>
<connection>
<GID>279</GID>
<name>IN_6</name></connection>
<intersection>-70.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>435 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-62,50,-62</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>455 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-97.5,50,-97.5</points>
<connection>
<GID>445</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>216 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8.5,1,-8.5,1.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>1.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-7.5,1.5,-7.5,2</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-8.5,1.5,-7.5,1.5</points>
<intersection>-8.5 0</intersection>
<intersection>-7.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>518 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-64,93.5,-64</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<connection>
<GID>326</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>218 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11.5,1.5,-11.5,2</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>1.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-10.5,1,-10.5,1.5</points>
<connection>
<GID>190</GID>
<name>IN_2</name></connection>
<intersection>1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-11.5,1.5,-10.5,1.5</points>
<intersection>-11.5 0</intersection>
<intersection>-10.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>276 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-62.5,7,-62</points>
<connection>
<GID>215</GID>
<name>IN_2</name></connection>
<intersection>-62 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>6.5,-62,6.5,-61.5</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>-62 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-62,7,-62</points>
<intersection>6.5 1</intersection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>243 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-40.5,8,-40</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>-40 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>9.5,-40,9.5,-39.5</points>
<connection>
<GID>173</GID>
<name>OUT_3</name></connection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>8,-40,9.5,-40</points>
<intersection>8 0</intersection>
<intersection>9.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>454 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-102.5,50,-102.5</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>457 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-100.5,50,-100.5</points>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>458 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-99.5,50,-99.5</points>
<connection>
<GID>460</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>456 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-98.5,50,-98.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>446 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-110.5,50,-110.5</points>
<connection>
<GID>455</GID>
<name>OUT_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>449 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-108.5,50,-108.5</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>450 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-107.5,50,-107.5</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>451 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-106,50,-106</points>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<intersection>50 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50,-106.5,50,-105.5</points>
<connection>
<GID>302</GID>
<name>IN_7</name></connection>
<connection>
<GID>302</GID>
<name>IN_6</name></connection>
<intersection>-106 1</intersection></vsegment></shape></wire>
<wire>
<ID>452 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-104.5,50,-104.5</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>453 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-103.5,50,-103.5</points>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>444 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>54.5,-95.5,54.5,-94.5</points>
<connection>
<GID>302</GID>
<name>SEL_0</name></connection>
<connection>
<GID>453</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>443 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-95.5,53.5,-89.5</points>
<connection>
<GID>302</GID>
<name>SEL_1</name></connection>
<connection>
<GID>238</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>441 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>52.5,-95.5,52.5,-94.5</points>
<connection>
<GID>302</GID>
<name>SEL_2</name></connection>
<connection>
<GID>454</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>442 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-95.5,51.5,-89.5</points>
<connection>
<GID>302</GID>
<name>SEL_3</name></connection>
<connection>
<GID>285</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>440 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56,-105,56.5,-105</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<connection>
<GID>395</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>380 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-110,-3,-105</points>
<connection>
<GID>235</GID>
<name>IN_1</name></connection>
<connection>
<GID>266</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>219 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,1,-13.5,2</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-13.5,1,-11.5,1</points>
<connection>
<GID>190</GID>
<name>IN_3</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>262 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>-1.5,-31.5,-1.5,-31</points>
<connection>
<GID>174</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>186</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>237 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-31.5,-9.5,-30.5</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<connection>
<GID>150</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>220 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-8,14,-7.5</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>12.5,-7.5,12.5,-7</points>
<connection>
<GID>189</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-7.5,14,-7.5</points>
<intersection>12.5 1</intersection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>374 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-110,-2,-110</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<connection>
<GID>415</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>221 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-7.5,11.5,-7</points>
<connection>
<GID>189</GID>
<name>OUT_1</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>12,-8,12,-7.5</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-7.5,12,-7.5</points>
<intersection>11.5 0</intersection>
<intersection>12 1</intersection></hsegment></shape></wire>
<wire>
<ID>524 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-95.5,98,-94.5</points>
<connection>
<GID>490</GID>
<name>SEL_0</name></connection>
<connection>
<GID>340</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>317 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-26,-43,-26</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<connection>
<GID>301</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>264 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>-3.5,-31.5,-3.5,-31</points>
<connection>
<GID>174</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>186</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>247 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-40.5,-9.5,-40</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>-40 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-8,-40,-8,-39.5</points>
<connection>
<GID>174</GID>
<name>OUT_3</name></connection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-9.5,-40,-8,-40</points>
<intersection>-9.5 0</intersection>
<intersection>-8 1</intersection></hsegment></shape></wire>
<wire>
<ID>222 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-7.5,10.5,-7</points>
<connection>
<GID>189</GID>
<name>OUT_2</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>10,-8,10,-7.5</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>10,-7.5,10.5,-7.5</points>
<intersection>10 1</intersection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>475 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,9.5,94.5,9.5</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<connection>
<GID>465</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>224 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-7.5,-5,-7</points>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-3.5,-8,-3.5,-7.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-5,-7.5,-3.5,-7.5</points>
<intersection>-5 0</intersection>
<intersection>-3.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>479 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,5.5,94.5,5.5</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<connection>
<GID>465</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>378 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-110,4,-105</points>
<connection>
<GID>235</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>418</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>225 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-8,-5.5,-7.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-6,-7.5,-6,-7</points>
<connection>
<GID>190</GID>
<name>OUT_1</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-6,-7.5,-5.5,-7.5</points>
<intersection>-6 1</intersection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>226 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-8,-7.5,-7.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-7,-7.5,-7,-7</points>
<connection>
<GID>190</GID>
<name>OUT_2</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-7.5,-7,-7.5</points>
<intersection>-7.5 0</intersection>
<intersection>-7 1</intersection></hsegment></shape></wire>
<wire>
<ID>318 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-24,-43,-24</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<connection>
<GID>301</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>260 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-1.5,-27,1.5,-27</points>
<connection>
<GID>186</GID>
<name>IN_3</name></connection>
<intersection>1.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1.5,-27,1.5,-25.5</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>-27 2</intersection></vsegment></shape></wire>
<wire>
<ID>227 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-8,-9.5,-7.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-8,-7.5,-8,-7</points>
<connection>
<GID>190</GID>
<name>OUT_3</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-9.5,-7.5,-8,-7.5</points>
<intersection>-9.5 0</intersection>
<intersection>-8 1</intersection></hsegment></shape></wire>
<wire>
<ID>322 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-36,-43,-36</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<connection>
<GID>336</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>228 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-2,20,-2</points>
<connection>
<GID>189</GID>
<name>carry_in</name></connection>
<intersection>20 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>20,-2.5,20,-2</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>-2 1</intersection></vsegment></shape></wire>
<wire>
<ID>382 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-110,-13.5,-110</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<connection>
<GID>401</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>229 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-8.5,-14.5,-4</points>
<connection>
<GID>190</GID>
<name>overflow</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-14.5,-8.5,-13,-8.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>230 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,-8.5,-15,-2</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15,-2,-14.5,-2</points>
<connection>
<GID>190</GID>
<name>carry_out</name></connection>
<intersection>-15 0</intersection></hsegment></shape></wire>
<wire>
<ID>236 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8.5,-31.5,-8.5,-31</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-7.5,-31,-7.5,-30.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-8.5,-31,-7.5,-31</points>
<intersection>-8.5 0</intersection>
<intersection>-7.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>325 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-40,-43,-40</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<connection>
<GID>319</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>238 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11.5,-31,-11.5,-30.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-10.5,-31.5,-10.5,-31</points>
<connection>
<GID>174</GID>
<name>IN_2</name></connection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-11.5,-31,-10.5,-31</points>
<intersection>-11.5 0</intersection>
<intersection>-10.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>240 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-40.5,14,-40</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>-40 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>12.5,-40,12.5,-39.5</points>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-40,14,-40</points>
<intersection>12.5 1</intersection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>320 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-34,-43,-34</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<connection>
<GID>333</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>366 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-91,-37,-91</points>
<connection>
<GID>381</GID>
<name>OUT</name></connection>
<connection>
<GID>392</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>213 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,1,-2.5,1.5</points>
<connection>
<GID>190</GID>
<name>IN_B_1</name></connection>
<intersection>1.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-0.5,1.5,-0.5,2</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-2.5,1.5,-0.5,1.5</points>
<intersection>-2.5 0</intersection>
<intersection>-0.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>266 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-34.5,20,-33.5</points>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-34.5,20,-34.5</points>
<connection>
<GID>173</GID>
<name>carry_in</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>241 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-40,11.5,-39.5</points>
<connection>
<GID>173</GID>
<name>OUT_1</name></connection>
<intersection>-40 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>12,-40.5,12,-40</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-40,12,-40</points>
<intersection>11.5 0</intersection>
<intersection>12 1</intersection></hsegment></shape></wire>
<wire>
<ID>242 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-40,10.5,-39.5</points>
<connection>
<GID>173</GID>
<name>OUT_2</name></connection>
<intersection>-40 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>10,-40.5,10,-40</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>10,-40,10.5,-40</points>
<intersection>10 1</intersection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>244 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-40,-5,-39.5</points>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection>
<intersection>-40 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-3.5,-40.5,-3.5,-40</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-5,-40,-3.5,-40</points>
<intersection>-5 0</intersection>
<intersection>-3.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>246 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-40.5,-7.5,-40</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>-40 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-7,-40,-7,-39.5</points>
<connection>
<GID>174</GID>
<name>OUT_2</name></connection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-40,-7,-40</points>
<intersection>-7.5 0</intersection>
<intersection>-7 1</intersection></hsegment></shape></wire>
<wire>
<ID>274 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-62.5,9,-62</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>-62 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>10.5,-62,10.5,-61.5</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>-62 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>9,-62,10.5,-62</points>
<intersection>9 0</intersection>
<intersection>10.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>249 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,-41,-15,-34.5</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15,-34.5,-14.5,-34.5</points>
<connection>
<GID>174</GID>
<name>carry_out</name></connection>
<intersection>-15 0</intersection></hsegment></shape></wire>
<wire>
<ID>232 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-31.5,9,-31</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>10.5,-31,10.5,-30.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>9,-31,10.5,-31</points>
<intersection>9 0</intersection>
<intersection>10.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>234 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-31.5,7,-31</points>
<connection>
<GID>173</GID>
<name>IN_2</name></connection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>6.5,-31,6.5,-30.5</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-31,7,-31</points>
<intersection>6.5 1</intersection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>278 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8.5,-62.5,-8.5,-62</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>-62 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-7.5,-62,-7.5,-61.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>-62 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-8.5,-62,-7.5,-62</points>
<intersection>-8.5 0</intersection>
<intersection>-7.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>253 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>16,-31.5,16,-31</points>
<connection>
<GID>173</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>183</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>284 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-16,-67.5,-14.5,-67.5</points>
<connection>
<GID>216</GID>
<name>overflow</name></connection>
<intersection>-16 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-16,-71.5,-16,-67.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>-67.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>251 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>15,-31.5,15,-31</points>
<connection>
<GID>173</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>183</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>252 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>14,-31.5,14,-31</points>
<connection>
<GID>173</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>183</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>250 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>13,-31.5,13,-31</points>
<connection>
<GID>173</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>376 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-110,3,-110</points>
<connection>
<GID>235</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>406</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>231 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1.5,-34.5,3,-34.5</points>
<connection>
<GID>174</GID>
<name>carry_in</name></connection>
<connection>
<GID>173</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>263 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>-2.5,-31.5,-2.5,-31</points>
<connection>
<GID>174</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>186</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>265 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>-4.5,-31.5,-4.5,-31</points>
<connection>
<GID>174</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>257 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-27,15,-26.5</points>
<connection>
<GID>183</GID>
<name>IN_2</name></connection>
<intersection>-26.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>17,-26.5,17,-25.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>15,-26.5,17,-26.5</points>
<intersection>15 0</intersection>
<intersection>17 1</intersection></hsegment></shape></wire>
<wire>
<ID>254 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-27,13,-25.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>362 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-75,-37,-75</points>
<connection>
<GID>376</GID>
<name>OUT</name></connection>
<connection>
<GID>385</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>209 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,1,8,1.5</points>
<connection>
<GID>189</GID>
<name>IN_1</name></connection>
<intersection>1.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>8.5,1.5,8.5,2</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>8,1.5,8.5,1.5</points>
<intersection>8 0</intersection>
<intersection>8.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>210 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,1,7,1.5</points>
<connection>
<GID>189</GID>
<name>IN_2</name></connection>
<intersection>1.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>6.5,1.5,6.5,2</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>6.5,1.5,7,1.5</points>
<intersection>6.5 1</intersection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>372 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-116,-8,-116</points>
<connection>
<GID>401</GID>
<name>in_A_less_B</name></connection>
<connection>
<GID>235</GID>
<name>A_less_B</name></connection></hsegment></shape></wire>
<wire>
<ID>211 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,1.5,4.5,2</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>1.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>6,1,6,1.5</points>
<connection>
<GID>189</GID>
<name>IN_3</name></connection>
<intersection>1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>4.5,1.5,6,1.5</points>
<intersection>4.5 0</intersection>
<intersection>6 1</intersection></hsegment></shape></wire>
<wire>
<ID>358 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-70,-43,-70</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<connection>
<GID>374</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>205 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,1,15,1.5</points>
<connection>
<GID>189</GID>
<name>IN_B_1</name></connection>
<intersection>1.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>17.5,1.5,17.5,2</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>15,1.5,17.5,1.5</points>
<intersection>15 0</intersection>
<intersection>17.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>529 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-108.5,93.5,-108.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>352 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-88,-43,-88</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<connection>
<GID>379</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>207 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>13,1,13,2</points>
<connection>
<GID>189</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>192</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>364 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-83,-37,-83</points>
<connection>
<GID>378</GID>
<name>OUT</name></connection>
<connection>
<GID>388</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>203 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1.5,-2,3,-2</points>
<connection>
<GID>190</GID>
<name>carry_in</name></connection>
<connection>
<GID>189</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>212 </ID>
<shape>
<vsegment>
<ID>1</ID>
<points>1.5,1,1.5,2</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,1,1.5,1</points>
<connection>
<GID>190</GID>
<name>IN_B_0</name></connection>
<intersection>1.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>513 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-68,93.5,-68</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<connection>
<GID>326</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>336 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-33,-37,-33</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<connection>
<GID>333</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>514 </ID>
<shape>
<hsegment>
<ID>7</ID>
<points>93,-67,93.5,-67</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<connection>
<GID>326</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>503 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>97,-60,97,-54</points>
<connection>
<GID>326</GID>
<name>SEL_1</name></connection>
<connection>
<GID>350</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>341 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-53,-37,-53</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<connection>
<GID>342</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>505 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-77,82.5,-56</points>
<intersection>-77 1</intersection>
<intersection>-76 4</intersection>
<intersection>-75 7</intersection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-77,93.5,-77</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>82.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72.5,-56,82.5,-56</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>82.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>82.5,-76,93.5,-76</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<intersection>82.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>82.5,-75,83.5,-75</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>349 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-80,-43,-80</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<connection>
<GID>377</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>517 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93,-65,93.5,-65</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<connection>
<GID>326</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>340 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-49,-37,-49</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<connection>
<GID>339</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>345 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-68,-43,-68</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<connection>
<GID>373</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>346 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-76,-43,-76</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<connection>
<GID>376</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>353 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-86,-43,-86</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<connection>
<GID>379</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>390 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,-117,-26.5,-116</points>
<connection>
<GID>401</GID>
<name>A_less_B</name></connection>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>-117 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-117,-26.5,-117</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<intersection>-26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>539 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-101.5,93.5,-101.5</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>279 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-62.5,-9.5,-61.5</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<connection>
<GID>208</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>348 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-78,-43,-78</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<connection>
<GID>377</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>525 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-112.5,82.5,-91.5</points>
<intersection>-112.5 1</intersection>
<intersection>-111.5 4</intersection>
<intersection>-110.5 7</intersection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-112.5,93.5,-112.5</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<intersection>82.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72.5,-91.5,82.5,-91.5</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>82.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>82.5,-111.5,93.5,-111.5</points>
<connection>
<GID>490</GID>
<name>IN_1</name></connection>
<intersection>82.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>82.5,-110.5,83.5,-110.5</points>
<connection>
<GID>491</GID>
<name>IN_0</name></connection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>280 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10.5,-62.5,-10.5,-61.5</points>
<connection>
<GID>216</GID>
<name>IN_2</name></connection>
<intersection>-61.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-11.5,-61.5,-10.5,-61.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>-10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>355 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-90,-43,-90</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<connection>
<GID>381</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>533 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-103.5,93.5,-103.5</points>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>356 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-96,-43,-96</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<connection>
<GID>382</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>281 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-62.5,-13.5,-61.5</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-13.5,-62.5,-11.5,-62.5</points>
<connection>
<GID>216</GID>
<name>IN_3</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>282 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>12.5,-81.5,12.5,-70.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<connection>
<GID>215</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>359 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-72,-43,-72</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<connection>
<GID>374</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>283 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-65.5,20,-65.5</points>
<connection>
<GID>213</GID>
<name>OUT_0</name></connection>
<connection>
<GID>215</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>357 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-94,-43,-94</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<connection>
<GID>382</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>275 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-62.5,8,-62</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>-62 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>8.5,-62,8.5,-61.5</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>-62 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>8,-62,8.5,-62</points>
<intersection>8 0</intersection>
<intersection>8.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>277 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-62,4.5,-61.5</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>-62 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>6,-62.5,6,-62</points>
<connection>
<GID>215</GID>
<name>IN_3</name></connection>
<intersection>-62 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-62,6,-62</points>
<intersection>4.5 0</intersection>
<intersection>6 1</intersection></hsegment></shape></wire>
<wire>
<ID>285 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>16,-62.5,17,-62.5</points>
<connection>
<GID>215</GID>
<name>IN_B_0</name></connection>
<intersection>17 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>17,-62.5,17,-61.5</points>
<connection>
<GID>220</GID>
<name>OUT_0</name></connection>
<intersection>-62.5 0</intersection></vsegment></shape></wire>
<wire>
<ID>287 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-62.5,13,-61.5</points>
<connection>
<GID>215</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>-62 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>13,-62,15,-62</points>
<intersection>13 0</intersection>
<intersection>14 5</intersection>
<intersection>15 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-62.5,15,-62</points>
<connection>
<GID>215</GID>
<name>IN_B_1</name></connection>
<intersection>-62 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>14,-62.5,14,-62</points>
<connection>
<GID>215</GID>
<name>IN_B_2</name></connection>
<intersection>-62 3</intersection></vsegment></shape></wire>
<wire>
<ID>288 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-70.5,11.5,-70.5</points>
<connection>
<GID>215</GID>
<name>OUT_1</name></connection>
<connection>
<GID>223</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>289 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-81.5,10.5,-70.5</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<connection>
<GID>215</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>290 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-70.5,9.5,-70.5</points>
<connection>
<GID>215</GID>
<name>OUT_3</name></connection>
<connection>
<GID>225</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>273 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1.5,-65.5,3,-65.5</points>
<connection>
<GID>216</GID>
<name>carry_in</name></connection>
<connection>
<GID>215</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>286 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,-62.5,-2.5,-61.5</points>
<connection>
<GID>216</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>-62 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-4.5,-62,-1.5,-62</points>
<intersection>-4.5 9</intersection>
<intersection>-3.5 10</intersection>
<intersection>-2.5 0</intersection>
<intersection>-1.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-1.5,-62.5,-1.5,-62</points>
<connection>
<GID>216</GID>
<name>IN_B_0</name></connection>
<intersection>-62 5</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-4.5,-62.5,-4.5,-62</points>
<connection>
<GID>216</GID>
<name>IN_B_3</name></connection>
<intersection>-62 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-3.5,-62.5,-3.5,-62</points>
<connection>
<GID>216</GID>
<name>IN_B_2</name></connection>
<intersection>-62 5</intersection></vsegment></shape></wire>
<wire>
<ID>291 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-70.5,-5,-70.5</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<connection>
<GID>226</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>292 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-81.5,-6,-70.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<connection>
<GID>216</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>293 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-70.5,-7,-70.5</points>
<connection>
<GID>216</GID>
<name>OUT_2</name></connection>
<connection>
<GID>228</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>294 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,-81.5,-8,-70.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<connection>
<GID>216</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>350 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-84,-43,-84</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<connection>
<GID>378</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>361 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-71,-37,-71</points>
<connection>
<GID>374</GID>
<name>OUT</name></connection>
<connection>
<GID>384</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>528 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-109.5,84,-93.5</points>
<intersection>-109.5 1</intersection>
<intersection>-93.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-109.5,88,-109.5</points>
<connection>
<GID>368</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72.5,-93.5,84,-93.5</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>490 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74,-35,94.5,-35</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<connection>
<GID>299</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>527 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>92,-109.5,93.5,-109.5</points>
<connection>
<GID>368</GID>
<name>OUT_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>351 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-82,-43,-82</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<connection>
<GID>361</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>386 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,-110,-20.5,-110</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<connection>
<GID>401</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>367 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-95,-37,-95</points>
<connection>
<GID>382</GID>
<name>OUT</name></connection>
<connection>
<GID>394</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>347 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-74,-43,-74</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>297 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,4,-43,4</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<connection>
<GID>232</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>296 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,2,-43,2</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<connection>
<GID>234</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>298 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,3,-37,3</points>
<connection>
<GID>231</GID>
<name>OUT</name></connection>
<connection>
<GID>236</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>408 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-37,41.5,-21</points>
<intersection>-37 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-37,45.5,-37</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-21,41.5,-21</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>516 </ID>
<shape>
<hsegment>
<ID>7</ID>
<points>93,-63,93.5,-63</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<connection>
<GID>326</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>309 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-12,-43,-12</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<connection>
<GID>271</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>308 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-14,-43,-14</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<connection>
<GID>274</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>310 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-13,-37,-13</points>
<connection>
<GID>268</GID>
<name>OUT</name></connection>
<connection>
<GID>275</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>375 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-110,-4,-110</points>
<connection>
<GID>235</GID>
<name>IN_2</name></connection>
<connection>
<GID>272</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>381 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-110,-5,-105</points>
<connection>
<GID>235</GID>
<name>IN_3</name></connection>
<connection>
<GID>419</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>379 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-110,2,-105</points>
<connection>
<GID>235</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>403</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>373 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-114,-8,-114</points>
<connection>
<GID>401</GID>
<name>in_A_equal_B</name></connection>
<connection>
<GID>235</GID>
<name>A_equal_B</name></connection></hsegment></shape></wire>
<wire>
<ID>371 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-112,-8,-112</points>
<connection>
<GID>401</GID>
<name>in_A_greater_B</name></connection>
<connection>
<GID>235</GID>
<name>A_greater_B</name></connection></hsegment></shape></wire>
<wire>
<ID>512 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>93,-69,93.5,-69</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<connection>
<GID>326</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>305 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-10,-43,-10</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<connection>
<GID>256</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>300 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,0,-43,0</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<connection>
<GID>240</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>299 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-2,-43,-2</points>
<connection>
<GID>237</GID>
<name>IN_1</name></connection>
<connection>
<GID>242</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>301 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-1,-37,-1</points>
<connection>
<GID>237</GID>
<name>OUT</name></connection>
<connection>
<GID>243</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>306 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-8,-43,-8</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<connection>
<GID>259</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>307 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-9,-37,-9</points>
<connection>
<GID>256</GID>
<name>OUT</name></connection>
<connection>
<GID>263</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>425 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-77,39,-56</points>
<intersection>-77 1</intersection>
<intersection>-76 4</intersection>
<intersection>-75 7</intersection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-77,50,-77</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-56,39,-56</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>39,-76,50,-76</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>39,-75,40,-75</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>426 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-75,50,-75</points>
<connection>
<GID>276</GID>
<name>OUT_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>409 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-36,51,-36</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>303 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-4,-43,-4</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<connection>
<GID>247</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>302 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-6,-43,-6</points>
<connection>
<GID>245</GID>
<name>IN_1</name></connection>
<connection>
<GID>250</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>304 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-5,-37,-5</points>
<connection>
<GID>245</GID>
<name>OUT</name></connection>
<connection>
<GID>251</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>509 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-73,93.5,-73</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<connection>
<GID>326</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>384 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-110,-14.5,-105</points>
<connection>
<GID>401</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>248</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>403 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-23,54.5,-17</points>
<connection>
<GID>433</GID>
<name>SEL_1</name></connection>
<connection>
<GID>249</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>385 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-110,-16.5,-105</points>
<connection>
<GID>401</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>284</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>412 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-32,51,-32</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>331 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-52,-43,-52</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<connection>
<GID>342</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>536 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>93,-98.5,93.5,-98.5</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>405 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-40,40,-19</points>
<intersection>-40 1</intersection>
<intersection>-39 4</intersection>
<intersection>-38 6</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-40,51,-40</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-19,40,-19</points>
<connection>
<GID>432</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>40,-39,51,-39</points>
<connection>
<GID>433</GID>
<name>IN_1</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>40,-38,41,-38</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>406 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-38,51,-38</points>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>462 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,11.5,96,17.5</points>
<connection>
<GID>465</GID>
<name>SEL_3</name></connection>
<connection>
<GID>257</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>411 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-33.5,51,-33.5</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>51 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>51,-34,51,-33</points>
<connection>
<GID>433</GID>
<name>IN_7</name></connection>
<connection>
<GID>433</GID>
<name>IN_6</name></connection>
<intersection>-33.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>464 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,11.5,99,12.5</points>
<connection>
<GID>465</GID>
<name>SEL_0</name></connection>
<connection>
<GID>265</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>469 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-1.5,94.5,-1.5</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<connection>
<GID>465</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>439 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-66,50,-66</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>434 </ID>
<shape>
<hsegment>
<ID>7</ID>
<points>49.5,-67,50,-67</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>438 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-64,50,-64</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>436 </ID>
<shape>
<hsegment>
<ID>7</ID>
<points>49.5,-63,50,-63</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>427 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-74,50,-74</points>
<connection>
<GID>448</GID>
<name>OUT_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>430 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-72,50,-72</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>433 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-68,50,-68</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>423 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-60,53.5,-54</points>
<connection>
<GID>279</GID>
<name>SEL_1</name></connection>
<connection>
<GID>446</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>422 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-60,51.5,-54</points>
<connection>
<GID>279</GID>
<name>SEL_3</name></connection>
<connection>
<GID>447</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>420 </ID>
<shape>
<hsegment>
<ID>7</ID>
<points>56,-69.5,56.5,-69.5</points>
<connection>
<GID>279</GID>
<name>OUT</name></connection>
<connection>
<GID>444</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>502 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>95,-60,95,-54</points>
<connection>
<GID>326</GID>
<name>SEL_3</name></connection>
<connection>
<GID>486</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>523 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-95.5,97,-89.5</points>
<connection>
<GID>490</GID>
<name>SEL_1</name></connection>
<connection>
<GID>281</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>468 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-2.5,85,13.5</points>
<intersection>-2.5 1</intersection>
<intersection>13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-2.5,89,-2.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,13.5,85,13.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>467 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>93,-2.5,94.5,-2.5</points>
<connection>
<GID>289</GID>
<name>OUT_0</name></connection>
<connection>
<GID>465</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>485 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-40,83.5,-19</points>
<intersection>-40 1</intersection>
<intersection>-39 4</intersection>
<intersection>-38 6</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-40,94.5,-40</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-19,83.5,-19</points>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>83.5,-39,94.5,-39</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>83.5,-38,84.5,-38</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>515 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-62,93.5,-62</points>
<connection>
<GID>489</GID>
<name>IN_0</name></connection>
<connection>
<GID>326</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>494 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-30,94.5,-30</points>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<connection>
<GID>299</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>499 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-29,94.5,-29</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<connection>
<GID>299</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>497 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-28,94.5,-28</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<connection>
<GID>299</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>535 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-97.5,93.5,-97.5</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>498 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-27,94.5,-27</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<connection>
<GID>299</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>496 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-26,94.5,-26</points>
<connection>
<GID>482</GID>
<name>IN_0</name></connection>
<connection>
<GID>299</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>495 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-25,94.5,-25</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<connection>
<GID>299</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>486 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88.5,-38,94.5,-38</points>
<connection>
<GID>412</GID>
<name>OUT_0</name></connection>
<connection>
<GID>299</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>487 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93,-37,94.5,-37</points>
<connection>
<GID>430</GID>
<name>OUT_0</name></connection>
<connection>
<GID>299</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>489 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-36,94.5,-36</points>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<connection>
<GID>299</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>491 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-33.5,94.5,-33.5</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<intersection>94.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>94.5,-34,94.5,-33</points>
<connection>
<GID>299</GID>
<name>IN_7</name></connection>
<connection>
<GID>299</GID>
<name>IN_6</name></connection>
<intersection>-33.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>492 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-32,94.5,-32</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<connection>
<GID>299</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>484 </ID>
<shape>
<vsegment>
<ID>4</ID>
<points>99,-23,99,-22</points>
<connection>
<GID>299</GID>
<name>SEL_0</name></connection>
<connection>
<GID>476</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>483 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>98,-23,98,-17</points>
<connection>
<GID>299</GID>
<name>SEL_1</name></connection>
<connection>
<GID>404</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>481 </ID>
<shape>
<vsegment>
<ID>4</ID>
<points>97,-23,97,-22</points>
<connection>
<GID>299</GID>
<name>SEL_2</name></connection>
<connection>
<GID>428</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>519 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-66,93.5,-66</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<connection>
<GID>326</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>482 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>96,-23,96,-17</points>
<connection>
<GID>299</GID>
<name>SEL_3</name></connection>
<connection>
<GID>477</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>319 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-25,-37,-25</points>
<connection>
<GID>301</GID>
<name>OUT</name></connection>
<connection>
<GID>307</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>477 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>94,6.5,94.5,6.5</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<connection>
<GID>465</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>328 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-48,-43,-48</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<connection>
<GID>339</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>321 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-32,-43,-32</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<connection>
<GID>333</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>488 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-37,85,-21</points>
<intersection>-37 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-37,89,-37</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-21,85,-21</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>323 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-38,-43,-38</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<connection>
<GID>336</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>332 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-56,-43,-56</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<connection>
<GID>322</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>324 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-42,-43,-42</points>
<connection>
<GID>319</GID>
<name>IN_1</name></connection>
<connection>
<GID>320</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>338 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-41,-37,-41</points>
<connection>
<GID>319</GID>
<name>OUT</name></connection>
<connection>
<GID>349</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>326 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-44,-43,-44</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<connection>
<GID>337</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>333 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-58,-43,-58</points>
<connection>
<GID>322</GID>
<name>IN_1</name></connection>
<connection>
<GID>329</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>342 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-57,-37,-57</points>
<connection>
<GID>322</GID>
<name>OUT</name></connection>
<connection>
<GID>355</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>327 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-46,-43,-46</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<connection>
<GID>337</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>329 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-50,-43,-50</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<connection>
<GID>339</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>506 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-75,93.5,-75</points>
<connection>
<GID>365</GID>
<name>OUT_0</name></connection>
<connection>
<GID>326</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>507 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>92,-74,93.5,-74</points>
<connection>
<GID>487</GID>
<name>OUT_0</name></connection>
<connection>
<GID>326</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>531 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-106,93.5,-106</points>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<intersection>93.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>93.5,-106.5,93.5,-105.5</points>
<connection>
<GID>490</GID>
<name>IN_7</name></connection>
<connection>
<GID>490</GID>
<name>IN_6</name></connection>
<intersection>-106 1</intersection></vsegment></shape></wire>
<wire>
<ID>510 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-72,93.5,-72</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<connection>
<GID>326</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>511 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-70.5,93.5,-70.5</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>93.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>93.5,-71,93.5,-70</points>
<connection>
<GID>326</GID>
<name>IN_7</name></connection>
<connection>
<GID>326</GID>
<name>IN_6</name></connection>
<intersection>-70.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>504 </ID>
<shape>
<vsegment>
<ID>4</ID>
<points>98,-60,98,-59</points>
<connection>
<GID>326</GID>
<name>SEL_0</name></connection>
<connection>
<GID>409</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>501 </ID>
<shape>
<vsegment>
<ID>4</ID>
<points>96,-60,96,-59</points>
<connection>
<GID>326</GID>
<name>SEL_2</name></connection>
<connection>
<GID>424</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>500 </ID>
<shape>
<hsegment>
<ID>9</ID>
<points>99.5,-69.5,100,-69.5</points>
<connection>
<GID>326</GID>
<name>OUT</name></connection>
<connection>
<GID>484</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>330 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-54,-43,-54</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<connection>
<GID>342</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>522 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-95.5,95,-89.5</points>
<connection>
<GID>490</GID>
<name>SEL_3</name></connection>
<connection>
<GID>328</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>335 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-62,-43,-62</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<connection>
<GID>343</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>337 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-37,-37,-37</points>
<connection>
<GID>336</GID>
<name>OUT</name></connection>
<connection>
<GID>348</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>339 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-45,-37,-45</points>
<connection>
<GID>337</GID>
<name>OUT</name></connection>
<connection>
<GID>351</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>343 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-61,-37,-61</points>
<connection>
<GID>343</GID>
<name>OUT</name></connection>
<connection>
<GID>357</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>363 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-79,-37,-79</points>
<connection>
<GID>377</GID>
<name>OUT</name></connection>
<connection>
<GID>386</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>365 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-87,-37,-87</points>
<connection>
<GID>379</GID>
<name>OUT</name></connection>
<connection>
<GID>391</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>391 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36.5,-114,-26.5,-114</points>
<connection>
<GID>401</GID>
<name>A_equal_B</name></connection>
<connection>
<GID>423</GID>
<name>IN_0</name></connection>
<intersection>-36.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-36.5,-115,-36.5,-113</points>
<connection>
<GID>425</GID>
<name>IN_1</name></connection>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<intersection>-114 1</intersection></vsegment></shape></wire>
<wire>
<ID>392 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,-112,-26.5,-111</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<connection>
<GID>401</GID>
<name>A_greater_B</name></connection>
<intersection>-111 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-111,-26.5,-111</points>
<connection>
<GID>393</GID>
<name>IN_1</name></connection>
<intersection>-26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>393 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-112,-42.5,-112</points>
<connection>
<GID>393</GID>
<name>OUT</name></connection>
<connection>
<GID>426</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>383 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-110,-15.5,-110</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<connection>
<GID>401</GID>
<name>IN_B_2</name></connection></vsegment></shape></wire>
<wire>
<ID>394 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-116,-42.5,-116</points>
<connection>
<GID>399</GID>
<name>IN_0</name></connection>
<connection>
<GID>425</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>389 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21.5,-110,-21.5,-105</points>
<connection>
<GID>401</GID>
<name>IN_1</name></connection>
<connection>
<GID>410</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>387 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-110,-22.5,-110</points>
<connection>
<GID>401</GID>
<name>IN_2</name></connection>
<connection>
<GID>407</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>388 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23.5,-110,-23.5,-105</points>
<connection>
<GID>401</GID>
<name>IN_3</name></connection>
<connection>
<GID>413</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>474 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>94,4.5,94.5,4.5</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<connection>
<GID>465</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>402 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-23,52.5,-17</points>
<connection>
<GID>433</GID>
<name>SEL_3</name></connection>
<connection>
<GID>414</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>400 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-32.5,57.5,-32.5</points>
<connection>
<GID>433</GID>
<name>OUT</name></connection>
<connection>
<GID>417</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>463 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,11.5,98,17.5</points>
<connection>
<GID>465</GID>
<name>SEL_1</name></connection>
<connection>
<GID>427</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>476 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>94,8.5,94.5,8.5</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<connection>
<GID>465</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>470 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74,-0.5,94.5,-0.5</points>
<connection>
<GID>431</GID>
<name>IN_0</name></connection>
<connection>
<GID>465</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>414 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-30,51,-30</points>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>419 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-29,51,-29</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>417 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-28,51,-28</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>418 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-27,51,-27</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>407 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-37,51,-37</points>
<connection>
<GID>437</GID>
<name>OUT_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>410 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-35,51,-35</points>
<connection>
<GID>438</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>413 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-31,51,-31</points>
<connection>
<GID>440</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>404 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>55.5,-23,55.5,-22</points>
<connection>
<GID>433</GID>
<name>SEL_0</name></connection>
<connection>
<GID>434</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>401 </ID>
<shape>
<vsegment>
<ID>2</ID>
<points>53.5,-23,53.5,-22</points>
<connection>
<GID>433</GID>
<name>SEL_2</name></connection>
<connection>
<GID>435</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>448 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-109.5,40.5,-93.5</points>
<intersection>-109.5 1</intersection>
<intersection>-93.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-109.5,44.5,-109.5</points>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-93.5,40.5,-93.5</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>465 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-5.5,83.5,15.5</points>
<intersection>-5.5 1</intersection>
<intersection>-4.5 4</intersection>
<intersection>-3.5 6</intersection>
<intersection>15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-5.5,94.5,-5.5</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,15.5,83.5,15.5</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>83.5,-4.5,94.5,-4.5</points>
<connection>
<GID>465</GID>
<name>IN_1</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>83.5,-3.5,84.5,-3.5</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>460 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>100.5,2,101,2</points>
<connection>
<GID>465</GID>
<name>OUT</name></connection>
<connection>
<GID>463</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>478 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,7.5,94.5,7.5</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<connection>
<GID>465</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>466 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88.5,-3.5,94.5,-3.5</points>
<connection>
<GID>468</GID>
<name>OUT_0</name></connection>
<connection>
<GID>465</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>471 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,1,94.5,1</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<intersection>94.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>94.5,0.5,94.5,1.5</points>
<connection>
<GID>465</GID>
<name>IN_7</name></connection>
<connection>
<GID>465</GID>
<name>IN_6</name></connection>
<intersection>1 1</intersection></vsegment></shape></wire>
<wire>
<ID>472 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>94,2.5,94.5,2.5</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<connection>
<GID>465</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>473 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,3.5,94.5,3.5</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<connection>
<GID>465</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>461 </ID>
<shape>
<vsegment>
<ID>4</ID>
<points>97,11.5,97,12.5</points>
<connection>
<GID>465</GID>
<name>SEL_2</name></connection>
<connection>
<GID>467</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>532 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>93,-104.5,93.5,-104.5</points>
<connection>
<GID>470</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>526 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-110.5,93.5,-110.5</points>
<connection>
<GID>491</GID>
<name>OUT_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_2</name></connection></hsegment></shape></wire></page 2></circuit>